magic
tech sky130A
magscale 1 2
timestamp 1712352531
<< nwell >>
rect -616 -797 616 797
<< mvpmos >>
rect -358 -500 -158 500
rect -100 -500 100 500
rect 158 -500 358 500
<< mvpdiff >>
rect -416 488 -358 500
rect -416 -488 -404 488
rect -370 -488 -358 488
rect -416 -500 -358 -488
rect -158 488 -100 500
rect -158 -488 -146 488
rect -112 -488 -100 488
rect -158 -500 -100 -488
rect 100 488 158 500
rect 100 -488 112 488
rect 146 -488 158 488
rect 100 -500 158 -488
rect 358 488 416 500
rect 358 -488 370 488
rect 404 -488 416 488
rect 358 -500 416 -488
<< mvpdiffc >>
rect -404 -488 -370 488
rect -146 -488 -112 488
rect 112 -488 146 488
rect 370 -488 404 488
<< mvnsubdiff >>
rect -550 719 550 731
rect -550 685 -442 719
rect 442 685 550 719
rect -550 673 550 685
rect -550 623 -492 673
rect -550 -623 -538 623
rect -504 -623 -492 623
rect 492 623 550 673
rect -550 -673 -492 -623
rect 492 -623 504 623
rect 538 -623 550 623
rect 492 -673 550 -623
rect -550 -685 550 -673
rect -550 -719 -442 -685
rect 442 -719 550 -685
rect -550 -731 550 -719
<< mvnsubdiffcont >>
rect -442 685 442 719
rect -538 -623 -504 623
rect 504 -623 538 623
rect -442 -719 442 -685
<< poly >>
rect -358 581 -158 597
rect -358 547 -342 581
rect -174 547 -158 581
rect -358 500 -158 547
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 500 100 547
rect 158 581 358 597
rect 158 547 174 581
rect 342 547 358 581
rect 158 500 358 547
rect -358 -547 -158 -500
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -358 -597 -158 -581
rect -100 -547 100 -500
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
rect 158 -547 358 -500
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 158 -597 358 -581
<< polycont >>
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
<< locali >>
rect -538 685 -442 719
rect 442 685 538 719
rect -538 623 -504 685
rect 504 623 538 685
rect -358 547 -342 581
rect -174 547 -158 581
rect -100 547 -84 581
rect 84 547 100 581
rect 158 547 174 581
rect 342 547 358 581
rect -404 488 -370 504
rect -404 -504 -370 -488
rect -146 488 -112 504
rect -146 -504 -112 -488
rect 112 488 146 504
rect 112 -504 146 -488
rect 370 488 404 504
rect 370 -504 404 -488
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect 158 -581 174 -547
rect 342 -581 358 -547
rect -538 -685 -504 -623
rect 504 -685 538 -623
rect -538 -719 -442 -685
rect 442 -719 538 -685
<< viali >>
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect -404 -488 -370 488
rect -146 -488 -112 488
rect 112 -488 146 488
rect 370 -488 404 488
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
<< metal1 >>
rect -354 581 -162 587
rect -354 547 -342 581
rect -174 547 -162 581
rect -354 541 -162 547
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect 162 581 354 587
rect 162 547 174 581
rect 342 547 354 581
rect 162 541 354 547
rect -410 488 -364 500
rect -410 -488 -404 488
rect -370 -488 -364 488
rect -410 -500 -364 -488
rect -152 488 -106 500
rect -152 -488 -146 488
rect -112 -488 -106 488
rect -152 -500 -106 -488
rect 106 488 152 500
rect 106 -488 112 488
rect 146 -488 152 488
rect 106 -500 152 -488
rect 364 488 410 500
rect 364 -488 370 488
rect 404 -488 410 488
rect 364 -500 410 -488
rect -354 -547 -162 -541
rect -354 -581 -342 -547
rect -174 -581 -162 -547
rect -354 -587 -162 -581
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
rect 162 -547 354 -541
rect 162 -581 174 -547
rect 342 -581 354 -547
rect 162 -587 354 -581
<< properties >>
string FIXED_BBOX -521 -702 521 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

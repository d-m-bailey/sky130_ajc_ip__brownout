magic
tech sky130A
magscale 1 2
timestamp 1712352531
<< nwell >>
rect -1119 -362 1119 362
<< mvpmos >>
rect -861 -136 -741 64
rect -683 -136 -563 64
rect -505 -136 -385 64
rect -327 -136 -207 64
rect -149 -136 -29 64
rect 29 -136 149 64
rect 207 -136 327 64
rect 385 -136 505 64
rect 563 -136 683 64
rect 741 -136 861 64
<< mvpdiff >>
rect -919 52 -861 64
rect -919 -124 -907 52
rect -873 -124 -861 52
rect -919 -136 -861 -124
rect -741 52 -683 64
rect -741 -124 -729 52
rect -695 -124 -683 52
rect -741 -136 -683 -124
rect -563 52 -505 64
rect -563 -124 -551 52
rect -517 -124 -505 52
rect -563 -136 -505 -124
rect -385 52 -327 64
rect -385 -124 -373 52
rect -339 -124 -327 52
rect -385 -136 -327 -124
rect -207 52 -149 64
rect -207 -124 -195 52
rect -161 -124 -149 52
rect -207 -136 -149 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 149 52 207 64
rect 149 -124 161 52
rect 195 -124 207 52
rect 149 -136 207 -124
rect 327 52 385 64
rect 327 -124 339 52
rect 373 -124 385 52
rect 327 -136 385 -124
rect 505 52 563 64
rect 505 -124 517 52
rect 551 -124 563 52
rect 505 -136 563 -124
rect 683 52 741 64
rect 683 -124 695 52
rect 729 -124 741 52
rect 683 -136 741 -124
rect 861 52 919 64
rect 861 -124 873 52
rect 907 -124 919 52
rect 861 -136 919 -124
<< mvpdiffc >>
rect -907 -124 -873 52
rect -729 -124 -695 52
rect -551 -124 -517 52
rect -373 -124 -339 52
rect -195 -124 -161 52
rect -17 -124 17 52
rect 161 -124 195 52
rect 339 -124 373 52
rect 517 -124 551 52
rect 695 -124 729 52
rect 873 -124 907 52
<< mvnsubdiff >>
rect -1053 284 1053 296
rect -1053 250 -945 284
rect 945 250 1053 284
rect -1053 238 1053 250
rect -1053 188 -995 238
rect -1053 -188 -1041 188
rect -1007 -188 -995 188
rect 995 188 1053 238
rect -1053 -238 -995 -188
rect 995 -188 1007 188
rect 1041 -188 1053 188
rect 995 -238 1053 -188
rect -1053 -250 1053 -238
rect -1053 -284 -945 -250
rect 945 -284 1053 -250
rect -1053 -296 1053 -284
<< mvnsubdiffcont >>
rect -945 250 945 284
rect -1041 -188 -1007 188
rect 1007 -188 1041 188
rect -945 -284 945 -250
<< poly >>
rect -861 145 -741 161
rect -861 111 -845 145
rect -757 111 -741 145
rect -861 64 -741 111
rect -683 145 -563 161
rect -683 111 -667 145
rect -579 111 -563 145
rect -683 64 -563 111
rect -505 145 -385 161
rect -505 111 -489 145
rect -401 111 -385 145
rect -505 64 -385 111
rect -327 145 -207 161
rect -327 111 -311 145
rect -223 111 -207 145
rect -327 64 -207 111
rect -149 145 -29 161
rect -149 111 -133 145
rect -45 111 -29 145
rect -149 64 -29 111
rect 29 145 149 161
rect 29 111 45 145
rect 133 111 149 145
rect 29 64 149 111
rect 207 145 327 161
rect 207 111 223 145
rect 311 111 327 145
rect 207 64 327 111
rect 385 145 505 161
rect 385 111 401 145
rect 489 111 505 145
rect 385 64 505 111
rect 563 145 683 161
rect 563 111 579 145
rect 667 111 683 145
rect 563 64 683 111
rect 741 145 861 161
rect 741 111 757 145
rect 845 111 861 145
rect 741 64 861 111
rect -861 -162 -741 -136
rect -683 -162 -563 -136
rect -505 -162 -385 -136
rect -327 -162 -207 -136
rect -149 -162 -29 -136
rect 29 -162 149 -136
rect 207 -162 327 -136
rect 385 -162 505 -136
rect 563 -162 683 -136
rect 741 -162 861 -136
<< polycont >>
rect -845 111 -757 145
rect -667 111 -579 145
rect -489 111 -401 145
rect -311 111 -223 145
rect -133 111 -45 145
rect 45 111 133 145
rect 223 111 311 145
rect 401 111 489 145
rect 579 111 667 145
rect 757 111 845 145
<< locali >>
rect -1041 250 -945 284
rect 945 250 1041 284
rect -1041 188 -1007 250
rect 1007 188 1041 250
rect -861 111 -845 145
rect -757 111 -741 145
rect -683 111 -667 145
rect -579 111 -563 145
rect -505 111 -489 145
rect -401 111 -385 145
rect -327 111 -311 145
rect -223 111 -207 145
rect -149 111 -133 145
rect -45 111 -29 145
rect 29 111 45 145
rect 133 111 149 145
rect 207 111 223 145
rect 311 111 327 145
rect 385 111 401 145
rect 489 111 505 145
rect 563 111 579 145
rect 667 111 683 145
rect 741 111 757 145
rect 845 111 861 145
rect -907 52 -873 68
rect -907 -140 -873 -124
rect -729 52 -695 68
rect -729 -140 -695 -124
rect -551 52 -517 68
rect -551 -140 -517 -124
rect -373 52 -339 68
rect -373 -140 -339 -124
rect -195 52 -161 68
rect -195 -140 -161 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 161 52 195 68
rect 161 -140 195 -124
rect 339 52 373 68
rect 339 -140 373 -124
rect 517 52 551 68
rect 517 -140 551 -124
rect 695 52 729 68
rect 695 -140 729 -124
rect 873 52 907 68
rect 873 -140 907 -124
rect -1041 -250 -1007 -188
rect 1007 -250 1041 -188
rect -1041 -284 -945 -250
rect 945 -284 1041 -250
<< viali >>
rect -845 111 -757 145
rect -667 111 -579 145
rect -489 111 -401 145
rect -311 111 -223 145
rect -133 111 -45 145
rect 45 111 133 145
rect 223 111 311 145
rect 401 111 489 145
rect 579 111 667 145
rect 757 111 845 145
rect -907 -124 -873 52
rect -729 -124 -695 52
rect -551 -124 -517 52
rect -373 -124 -339 52
rect -195 -124 -161 52
rect -17 -124 17 52
rect 161 -124 195 52
rect 339 -124 373 52
rect 517 -124 551 52
rect 695 -124 729 52
rect 873 -124 907 52
<< metal1 >>
rect -857 145 -745 151
rect -857 111 -845 145
rect -757 111 -745 145
rect -857 105 -745 111
rect -679 145 -567 151
rect -679 111 -667 145
rect -579 111 -567 145
rect -679 105 -567 111
rect -501 145 -389 151
rect -501 111 -489 145
rect -401 111 -389 145
rect -501 105 -389 111
rect -323 145 -211 151
rect -323 111 -311 145
rect -223 111 -211 145
rect -323 105 -211 111
rect -145 145 -33 151
rect -145 111 -133 145
rect -45 111 -33 145
rect -145 105 -33 111
rect 33 145 145 151
rect 33 111 45 145
rect 133 111 145 145
rect 33 105 145 111
rect 211 145 323 151
rect 211 111 223 145
rect 311 111 323 145
rect 211 105 323 111
rect 389 145 501 151
rect 389 111 401 145
rect 489 111 501 145
rect 389 105 501 111
rect 567 145 679 151
rect 567 111 579 145
rect 667 111 679 145
rect 567 105 679 111
rect 745 145 857 151
rect 745 111 757 145
rect 845 111 857 145
rect 745 105 857 111
rect -913 52 -867 64
rect -913 -124 -907 52
rect -873 -124 -867 52
rect -913 -136 -867 -124
rect -735 52 -689 64
rect -735 -124 -729 52
rect -695 -124 -689 52
rect -735 -136 -689 -124
rect -557 52 -511 64
rect -557 -124 -551 52
rect -517 -124 -511 52
rect -557 -136 -511 -124
rect -379 52 -333 64
rect -379 -124 -373 52
rect -339 -124 -333 52
rect -379 -136 -333 -124
rect -201 52 -155 64
rect -201 -124 -195 52
rect -161 -124 -155 52
rect -201 -136 -155 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 155 52 201 64
rect 155 -124 161 52
rect 195 -124 201 52
rect 155 -136 201 -124
rect 333 52 379 64
rect 333 -124 339 52
rect 373 -124 379 52
rect 333 -136 379 -124
rect 511 52 557 64
rect 511 -124 517 52
rect 551 -124 557 52
rect 511 -136 557 -124
rect 689 52 735 64
rect 689 -124 695 52
rect 729 -124 735 52
rect 689 -136 735 -124
rect 867 52 913 64
rect 867 -124 873 52
rect 907 -124 913 52
rect 867 -136 913 -124
<< properties >>
string FIXED_BBOX -1024 -267 1024 267
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.6 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

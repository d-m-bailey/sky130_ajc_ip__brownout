magic
tech sky130A
magscale 1 2
timestamp 1712352531
<< pwell >>
rect -5173 -1109 5173 1109
<< mvnmos >>
rect -4945 767 -3345 851
rect -3287 767 -1687 851
rect -1629 767 -29 851
rect 29 767 1629 851
rect 1687 767 3287 851
rect 3345 767 4945 851
rect -4945 527 -3345 611
rect -3287 527 -1687 611
rect -1629 527 -29 611
rect 29 527 1629 611
rect 1687 527 3287 611
rect 3345 527 4945 611
rect -4945 287 -3345 371
rect -3287 287 -1687 371
rect -1629 287 -29 371
rect 29 287 1629 371
rect 1687 287 3287 371
rect 3345 287 4945 371
rect -4945 47 -3345 131
rect -3287 47 -1687 131
rect -1629 47 -29 131
rect 29 47 1629 131
rect 1687 47 3287 131
rect 3345 47 4945 131
rect -4945 -193 -3345 -109
rect -3287 -193 -1687 -109
rect -1629 -193 -29 -109
rect 29 -193 1629 -109
rect 1687 -193 3287 -109
rect 3345 -193 4945 -109
rect -4945 -433 -3345 -349
rect -3287 -433 -1687 -349
rect -1629 -433 -29 -349
rect 29 -433 1629 -349
rect 1687 -433 3287 -349
rect 3345 -433 4945 -349
rect -4945 -673 -3345 -589
rect -3287 -673 -1687 -589
rect -1629 -673 -29 -589
rect 29 -673 1629 -589
rect 1687 -673 3287 -589
rect 3345 -673 4945 -589
rect -4945 -913 -3345 -829
rect -3287 -913 -1687 -829
rect -1629 -913 -29 -829
rect 29 -913 1629 -829
rect 1687 -913 3287 -829
rect 3345 -913 4945 -829
<< mvndiff >>
rect -5003 839 -4945 851
rect -5003 779 -4991 839
rect -4957 779 -4945 839
rect -5003 767 -4945 779
rect -3345 839 -3287 851
rect -3345 779 -3333 839
rect -3299 779 -3287 839
rect -3345 767 -3287 779
rect -1687 839 -1629 851
rect -1687 779 -1675 839
rect -1641 779 -1629 839
rect -1687 767 -1629 779
rect -29 839 29 851
rect -29 779 -17 839
rect 17 779 29 839
rect -29 767 29 779
rect 1629 839 1687 851
rect 1629 779 1641 839
rect 1675 779 1687 839
rect 1629 767 1687 779
rect 3287 839 3345 851
rect 3287 779 3299 839
rect 3333 779 3345 839
rect 3287 767 3345 779
rect 4945 839 5003 851
rect 4945 779 4957 839
rect 4991 779 5003 839
rect 4945 767 5003 779
rect -5003 599 -4945 611
rect -5003 539 -4991 599
rect -4957 539 -4945 599
rect -5003 527 -4945 539
rect -3345 599 -3287 611
rect -3345 539 -3333 599
rect -3299 539 -3287 599
rect -3345 527 -3287 539
rect -1687 599 -1629 611
rect -1687 539 -1675 599
rect -1641 539 -1629 599
rect -1687 527 -1629 539
rect -29 599 29 611
rect -29 539 -17 599
rect 17 539 29 599
rect -29 527 29 539
rect 1629 599 1687 611
rect 1629 539 1641 599
rect 1675 539 1687 599
rect 1629 527 1687 539
rect 3287 599 3345 611
rect 3287 539 3299 599
rect 3333 539 3345 599
rect 3287 527 3345 539
rect 4945 599 5003 611
rect 4945 539 4957 599
rect 4991 539 5003 599
rect 4945 527 5003 539
rect -5003 359 -4945 371
rect -5003 299 -4991 359
rect -4957 299 -4945 359
rect -5003 287 -4945 299
rect -3345 359 -3287 371
rect -3345 299 -3333 359
rect -3299 299 -3287 359
rect -3345 287 -3287 299
rect -1687 359 -1629 371
rect -1687 299 -1675 359
rect -1641 299 -1629 359
rect -1687 287 -1629 299
rect -29 359 29 371
rect -29 299 -17 359
rect 17 299 29 359
rect -29 287 29 299
rect 1629 359 1687 371
rect 1629 299 1641 359
rect 1675 299 1687 359
rect 1629 287 1687 299
rect 3287 359 3345 371
rect 3287 299 3299 359
rect 3333 299 3345 359
rect 3287 287 3345 299
rect 4945 359 5003 371
rect 4945 299 4957 359
rect 4991 299 5003 359
rect 4945 287 5003 299
rect -5003 119 -4945 131
rect -5003 59 -4991 119
rect -4957 59 -4945 119
rect -5003 47 -4945 59
rect -3345 119 -3287 131
rect -3345 59 -3333 119
rect -3299 59 -3287 119
rect -3345 47 -3287 59
rect -1687 119 -1629 131
rect -1687 59 -1675 119
rect -1641 59 -1629 119
rect -1687 47 -1629 59
rect -29 119 29 131
rect -29 59 -17 119
rect 17 59 29 119
rect -29 47 29 59
rect 1629 119 1687 131
rect 1629 59 1641 119
rect 1675 59 1687 119
rect 1629 47 1687 59
rect 3287 119 3345 131
rect 3287 59 3299 119
rect 3333 59 3345 119
rect 3287 47 3345 59
rect 4945 119 5003 131
rect 4945 59 4957 119
rect 4991 59 5003 119
rect 4945 47 5003 59
rect -5003 -121 -4945 -109
rect -5003 -181 -4991 -121
rect -4957 -181 -4945 -121
rect -5003 -193 -4945 -181
rect -3345 -121 -3287 -109
rect -3345 -181 -3333 -121
rect -3299 -181 -3287 -121
rect -3345 -193 -3287 -181
rect -1687 -121 -1629 -109
rect -1687 -181 -1675 -121
rect -1641 -181 -1629 -121
rect -1687 -193 -1629 -181
rect -29 -121 29 -109
rect -29 -181 -17 -121
rect 17 -181 29 -121
rect -29 -193 29 -181
rect 1629 -121 1687 -109
rect 1629 -181 1641 -121
rect 1675 -181 1687 -121
rect 1629 -193 1687 -181
rect 3287 -121 3345 -109
rect 3287 -181 3299 -121
rect 3333 -181 3345 -121
rect 3287 -193 3345 -181
rect 4945 -121 5003 -109
rect 4945 -181 4957 -121
rect 4991 -181 5003 -121
rect 4945 -193 5003 -181
rect -5003 -361 -4945 -349
rect -5003 -421 -4991 -361
rect -4957 -421 -4945 -361
rect -5003 -433 -4945 -421
rect -3345 -361 -3287 -349
rect -3345 -421 -3333 -361
rect -3299 -421 -3287 -361
rect -3345 -433 -3287 -421
rect -1687 -361 -1629 -349
rect -1687 -421 -1675 -361
rect -1641 -421 -1629 -361
rect -1687 -433 -1629 -421
rect -29 -361 29 -349
rect -29 -421 -17 -361
rect 17 -421 29 -361
rect -29 -433 29 -421
rect 1629 -361 1687 -349
rect 1629 -421 1641 -361
rect 1675 -421 1687 -361
rect 1629 -433 1687 -421
rect 3287 -361 3345 -349
rect 3287 -421 3299 -361
rect 3333 -421 3345 -361
rect 3287 -433 3345 -421
rect 4945 -361 5003 -349
rect 4945 -421 4957 -361
rect 4991 -421 5003 -361
rect 4945 -433 5003 -421
rect -5003 -601 -4945 -589
rect -5003 -661 -4991 -601
rect -4957 -661 -4945 -601
rect -5003 -673 -4945 -661
rect -3345 -601 -3287 -589
rect -3345 -661 -3333 -601
rect -3299 -661 -3287 -601
rect -3345 -673 -3287 -661
rect -1687 -601 -1629 -589
rect -1687 -661 -1675 -601
rect -1641 -661 -1629 -601
rect -1687 -673 -1629 -661
rect -29 -601 29 -589
rect -29 -661 -17 -601
rect 17 -661 29 -601
rect -29 -673 29 -661
rect 1629 -601 1687 -589
rect 1629 -661 1641 -601
rect 1675 -661 1687 -601
rect 1629 -673 1687 -661
rect 3287 -601 3345 -589
rect 3287 -661 3299 -601
rect 3333 -661 3345 -601
rect 3287 -673 3345 -661
rect 4945 -601 5003 -589
rect 4945 -661 4957 -601
rect 4991 -661 5003 -601
rect 4945 -673 5003 -661
rect -5003 -841 -4945 -829
rect -5003 -901 -4991 -841
rect -4957 -901 -4945 -841
rect -5003 -913 -4945 -901
rect -3345 -841 -3287 -829
rect -3345 -901 -3333 -841
rect -3299 -901 -3287 -841
rect -3345 -913 -3287 -901
rect -1687 -841 -1629 -829
rect -1687 -901 -1675 -841
rect -1641 -901 -1629 -841
rect -1687 -913 -1629 -901
rect -29 -841 29 -829
rect -29 -901 -17 -841
rect 17 -901 29 -841
rect -29 -913 29 -901
rect 1629 -841 1687 -829
rect 1629 -901 1641 -841
rect 1675 -901 1687 -841
rect 1629 -913 1687 -901
rect 3287 -841 3345 -829
rect 3287 -901 3299 -841
rect 3333 -901 3345 -841
rect 3287 -913 3345 -901
rect 4945 -841 5003 -829
rect 4945 -901 4957 -841
rect 4991 -901 5003 -841
rect 4945 -913 5003 -901
<< mvndiffc >>
rect -4991 779 -4957 839
rect -3333 779 -3299 839
rect -1675 779 -1641 839
rect -17 779 17 839
rect 1641 779 1675 839
rect 3299 779 3333 839
rect 4957 779 4991 839
rect -4991 539 -4957 599
rect -3333 539 -3299 599
rect -1675 539 -1641 599
rect -17 539 17 599
rect 1641 539 1675 599
rect 3299 539 3333 599
rect 4957 539 4991 599
rect -4991 299 -4957 359
rect -3333 299 -3299 359
rect -1675 299 -1641 359
rect -17 299 17 359
rect 1641 299 1675 359
rect 3299 299 3333 359
rect 4957 299 4991 359
rect -4991 59 -4957 119
rect -3333 59 -3299 119
rect -1675 59 -1641 119
rect -17 59 17 119
rect 1641 59 1675 119
rect 3299 59 3333 119
rect 4957 59 4991 119
rect -4991 -181 -4957 -121
rect -3333 -181 -3299 -121
rect -1675 -181 -1641 -121
rect -17 -181 17 -121
rect 1641 -181 1675 -121
rect 3299 -181 3333 -121
rect 4957 -181 4991 -121
rect -4991 -421 -4957 -361
rect -3333 -421 -3299 -361
rect -1675 -421 -1641 -361
rect -17 -421 17 -361
rect 1641 -421 1675 -361
rect 3299 -421 3333 -361
rect 4957 -421 4991 -361
rect -4991 -661 -4957 -601
rect -3333 -661 -3299 -601
rect -1675 -661 -1641 -601
rect -17 -661 17 -601
rect 1641 -661 1675 -601
rect 3299 -661 3333 -601
rect 4957 -661 4991 -601
rect -4991 -901 -4957 -841
rect -3333 -901 -3299 -841
rect -1675 -901 -1641 -841
rect -17 -901 17 -841
rect 1641 -901 1675 -841
rect 3299 -901 3333 -841
rect 4957 -901 4991 -841
<< mvpsubdiff >>
rect -5137 1061 5137 1073
rect -5137 1027 -5029 1061
rect 5029 1027 5137 1061
rect -5137 1015 5137 1027
rect -5137 965 -5079 1015
rect -5137 -965 -5125 965
rect -5091 -965 -5079 965
rect 5079 965 5137 1015
rect -5137 -1015 -5079 -965
rect 5079 -965 5091 965
rect 5125 -965 5137 965
rect 5079 -1015 5137 -965
rect -5137 -1027 5137 -1015
rect -5137 -1061 -5029 -1027
rect 5029 -1061 5137 -1027
rect -5137 -1073 5137 -1061
<< mvpsubdiffcont >>
rect -5029 1027 5029 1061
rect -5125 -965 -5091 965
rect 5091 -965 5125 965
rect -5029 -1061 5029 -1027
<< poly >>
rect -4945 923 -3345 939
rect -4945 889 -4929 923
rect -3361 889 -3345 923
rect -4945 851 -3345 889
rect -3287 923 -1687 939
rect -3287 889 -3271 923
rect -1703 889 -1687 923
rect -3287 851 -1687 889
rect -1629 923 -29 939
rect -1629 889 -1613 923
rect -45 889 -29 923
rect -1629 851 -29 889
rect 29 923 1629 939
rect 29 889 45 923
rect 1613 889 1629 923
rect 29 851 1629 889
rect 1687 923 3287 939
rect 1687 889 1703 923
rect 3271 889 3287 923
rect 1687 851 3287 889
rect 3345 923 4945 939
rect 3345 889 3361 923
rect 4929 889 4945 923
rect 3345 851 4945 889
rect -4945 741 -3345 767
rect -3287 741 -1687 767
rect -1629 741 -29 767
rect 29 741 1629 767
rect 1687 741 3287 767
rect 3345 741 4945 767
rect -4945 683 -3345 699
rect -4945 649 -4929 683
rect -3361 649 -3345 683
rect -4945 611 -3345 649
rect -3287 683 -1687 699
rect -3287 649 -3271 683
rect -1703 649 -1687 683
rect -3287 611 -1687 649
rect -1629 683 -29 699
rect -1629 649 -1613 683
rect -45 649 -29 683
rect -1629 611 -29 649
rect 29 683 1629 699
rect 29 649 45 683
rect 1613 649 1629 683
rect 29 611 1629 649
rect 1687 683 3287 699
rect 1687 649 1703 683
rect 3271 649 3287 683
rect 1687 611 3287 649
rect 3345 683 4945 699
rect 3345 649 3361 683
rect 4929 649 4945 683
rect 3345 611 4945 649
rect -4945 501 -3345 527
rect -3287 501 -1687 527
rect -1629 501 -29 527
rect 29 501 1629 527
rect 1687 501 3287 527
rect 3345 501 4945 527
rect -4945 443 -3345 459
rect -4945 409 -4929 443
rect -3361 409 -3345 443
rect -4945 371 -3345 409
rect -3287 443 -1687 459
rect -3287 409 -3271 443
rect -1703 409 -1687 443
rect -3287 371 -1687 409
rect -1629 443 -29 459
rect -1629 409 -1613 443
rect -45 409 -29 443
rect -1629 371 -29 409
rect 29 443 1629 459
rect 29 409 45 443
rect 1613 409 1629 443
rect 29 371 1629 409
rect 1687 443 3287 459
rect 1687 409 1703 443
rect 3271 409 3287 443
rect 1687 371 3287 409
rect 3345 443 4945 459
rect 3345 409 3361 443
rect 4929 409 4945 443
rect 3345 371 4945 409
rect -4945 261 -3345 287
rect -3287 261 -1687 287
rect -1629 261 -29 287
rect 29 261 1629 287
rect 1687 261 3287 287
rect 3345 261 4945 287
rect -4945 203 -3345 219
rect -4945 169 -4929 203
rect -3361 169 -3345 203
rect -4945 131 -3345 169
rect -3287 203 -1687 219
rect -3287 169 -3271 203
rect -1703 169 -1687 203
rect -3287 131 -1687 169
rect -1629 203 -29 219
rect -1629 169 -1613 203
rect -45 169 -29 203
rect -1629 131 -29 169
rect 29 203 1629 219
rect 29 169 45 203
rect 1613 169 1629 203
rect 29 131 1629 169
rect 1687 203 3287 219
rect 1687 169 1703 203
rect 3271 169 3287 203
rect 1687 131 3287 169
rect 3345 203 4945 219
rect 3345 169 3361 203
rect 4929 169 4945 203
rect 3345 131 4945 169
rect -4945 21 -3345 47
rect -3287 21 -1687 47
rect -1629 21 -29 47
rect 29 21 1629 47
rect 1687 21 3287 47
rect 3345 21 4945 47
rect -4945 -37 -3345 -21
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -4945 -109 -3345 -71
rect -3287 -37 -1687 -21
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -3287 -109 -1687 -71
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -109 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -109 1629 -71
rect 1687 -37 3287 -21
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 1687 -109 3287 -71
rect 3345 -37 4945 -21
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 3345 -109 4945 -71
rect -4945 -219 -3345 -193
rect -3287 -219 -1687 -193
rect -1629 -219 -29 -193
rect 29 -219 1629 -193
rect 1687 -219 3287 -193
rect 3345 -219 4945 -193
rect -4945 -277 -3345 -261
rect -4945 -311 -4929 -277
rect -3361 -311 -3345 -277
rect -4945 -349 -3345 -311
rect -3287 -277 -1687 -261
rect -3287 -311 -3271 -277
rect -1703 -311 -1687 -277
rect -3287 -349 -1687 -311
rect -1629 -277 -29 -261
rect -1629 -311 -1613 -277
rect -45 -311 -29 -277
rect -1629 -349 -29 -311
rect 29 -277 1629 -261
rect 29 -311 45 -277
rect 1613 -311 1629 -277
rect 29 -349 1629 -311
rect 1687 -277 3287 -261
rect 1687 -311 1703 -277
rect 3271 -311 3287 -277
rect 1687 -349 3287 -311
rect 3345 -277 4945 -261
rect 3345 -311 3361 -277
rect 4929 -311 4945 -277
rect 3345 -349 4945 -311
rect -4945 -459 -3345 -433
rect -3287 -459 -1687 -433
rect -1629 -459 -29 -433
rect 29 -459 1629 -433
rect 1687 -459 3287 -433
rect 3345 -459 4945 -433
rect -4945 -517 -3345 -501
rect -4945 -551 -4929 -517
rect -3361 -551 -3345 -517
rect -4945 -589 -3345 -551
rect -3287 -517 -1687 -501
rect -3287 -551 -3271 -517
rect -1703 -551 -1687 -517
rect -3287 -589 -1687 -551
rect -1629 -517 -29 -501
rect -1629 -551 -1613 -517
rect -45 -551 -29 -517
rect -1629 -589 -29 -551
rect 29 -517 1629 -501
rect 29 -551 45 -517
rect 1613 -551 1629 -517
rect 29 -589 1629 -551
rect 1687 -517 3287 -501
rect 1687 -551 1703 -517
rect 3271 -551 3287 -517
rect 1687 -589 3287 -551
rect 3345 -517 4945 -501
rect 3345 -551 3361 -517
rect 4929 -551 4945 -517
rect 3345 -589 4945 -551
rect -4945 -699 -3345 -673
rect -3287 -699 -1687 -673
rect -1629 -699 -29 -673
rect 29 -699 1629 -673
rect 1687 -699 3287 -673
rect 3345 -699 4945 -673
rect -4945 -757 -3345 -741
rect -4945 -791 -4929 -757
rect -3361 -791 -3345 -757
rect -4945 -829 -3345 -791
rect -3287 -757 -1687 -741
rect -3287 -791 -3271 -757
rect -1703 -791 -1687 -757
rect -3287 -829 -1687 -791
rect -1629 -757 -29 -741
rect -1629 -791 -1613 -757
rect -45 -791 -29 -757
rect -1629 -829 -29 -791
rect 29 -757 1629 -741
rect 29 -791 45 -757
rect 1613 -791 1629 -757
rect 29 -829 1629 -791
rect 1687 -757 3287 -741
rect 1687 -791 1703 -757
rect 3271 -791 3287 -757
rect 1687 -829 3287 -791
rect 3345 -757 4945 -741
rect 3345 -791 3361 -757
rect 4929 -791 4945 -757
rect 3345 -829 4945 -791
rect -4945 -939 -3345 -913
rect -3287 -939 -1687 -913
rect -1629 -939 -29 -913
rect 29 -939 1629 -913
rect 1687 -939 3287 -913
rect 3345 -939 4945 -913
<< polycont >>
rect -4929 889 -3361 923
rect -3271 889 -1703 923
rect -1613 889 -45 923
rect 45 889 1613 923
rect 1703 889 3271 923
rect 3361 889 4929 923
rect -4929 649 -3361 683
rect -3271 649 -1703 683
rect -1613 649 -45 683
rect 45 649 1613 683
rect 1703 649 3271 683
rect 3361 649 4929 683
rect -4929 409 -3361 443
rect -3271 409 -1703 443
rect -1613 409 -45 443
rect 45 409 1613 443
rect 1703 409 3271 443
rect 3361 409 4929 443
rect -4929 169 -3361 203
rect -3271 169 -1703 203
rect -1613 169 -45 203
rect 45 169 1613 203
rect 1703 169 3271 203
rect 3361 169 4929 203
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect -4929 -311 -3361 -277
rect -3271 -311 -1703 -277
rect -1613 -311 -45 -277
rect 45 -311 1613 -277
rect 1703 -311 3271 -277
rect 3361 -311 4929 -277
rect -4929 -551 -3361 -517
rect -3271 -551 -1703 -517
rect -1613 -551 -45 -517
rect 45 -551 1613 -517
rect 1703 -551 3271 -517
rect 3361 -551 4929 -517
rect -4929 -791 -3361 -757
rect -3271 -791 -1703 -757
rect -1613 -791 -45 -757
rect 45 -791 1613 -757
rect 1703 -791 3271 -757
rect 3361 -791 4929 -757
<< locali >>
rect -5125 1027 -5029 1061
rect 5029 1027 5125 1061
rect -5125 965 -5091 1027
rect 5091 965 5125 1027
rect -4945 889 -4929 923
rect -3361 889 -3345 923
rect -3287 889 -3271 923
rect -1703 889 -1687 923
rect -1629 889 -1613 923
rect -45 889 -29 923
rect 29 889 45 923
rect 1613 889 1629 923
rect 1687 889 1703 923
rect 3271 889 3287 923
rect 3345 889 3361 923
rect 4929 889 4945 923
rect -4991 839 -4957 855
rect -4991 763 -4957 779
rect -3333 839 -3299 855
rect -3333 763 -3299 779
rect -1675 839 -1641 855
rect -1675 763 -1641 779
rect -17 839 17 855
rect -17 763 17 779
rect 1641 839 1675 855
rect 1641 763 1675 779
rect 3299 839 3333 855
rect 3299 763 3333 779
rect 4957 839 4991 855
rect 4957 763 4991 779
rect -4945 649 -4929 683
rect -3361 649 -3345 683
rect -3287 649 -3271 683
rect -1703 649 -1687 683
rect -1629 649 -1613 683
rect -45 649 -29 683
rect 29 649 45 683
rect 1613 649 1629 683
rect 1687 649 1703 683
rect 3271 649 3287 683
rect 3345 649 3361 683
rect 4929 649 4945 683
rect -4991 599 -4957 615
rect -4991 523 -4957 539
rect -3333 599 -3299 615
rect -3333 523 -3299 539
rect -1675 599 -1641 615
rect -1675 523 -1641 539
rect -17 599 17 615
rect -17 523 17 539
rect 1641 599 1675 615
rect 1641 523 1675 539
rect 3299 599 3333 615
rect 3299 523 3333 539
rect 4957 599 4991 615
rect 4957 523 4991 539
rect -4945 409 -4929 443
rect -3361 409 -3345 443
rect -3287 409 -3271 443
rect -1703 409 -1687 443
rect -1629 409 -1613 443
rect -45 409 -29 443
rect 29 409 45 443
rect 1613 409 1629 443
rect 1687 409 1703 443
rect 3271 409 3287 443
rect 3345 409 3361 443
rect 4929 409 4945 443
rect -4991 359 -4957 375
rect -4991 283 -4957 299
rect -3333 359 -3299 375
rect -3333 283 -3299 299
rect -1675 359 -1641 375
rect -1675 283 -1641 299
rect -17 359 17 375
rect -17 283 17 299
rect 1641 359 1675 375
rect 1641 283 1675 299
rect 3299 359 3333 375
rect 3299 283 3333 299
rect 4957 359 4991 375
rect 4957 283 4991 299
rect -4945 169 -4929 203
rect -3361 169 -3345 203
rect -3287 169 -3271 203
rect -1703 169 -1687 203
rect -1629 169 -1613 203
rect -45 169 -29 203
rect 29 169 45 203
rect 1613 169 1629 203
rect 1687 169 1703 203
rect 3271 169 3287 203
rect 3345 169 3361 203
rect 4929 169 4945 203
rect -4991 119 -4957 135
rect -4991 43 -4957 59
rect -3333 119 -3299 135
rect -3333 43 -3299 59
rect -1675 119 -1641 135
rect -1675 43 -1641 59
rect -17 119 17 135
rect -17 43 17 59
rect 1641 119 1675 135
rect 1641 43 1675 59
rect 3299 119 3333 135
rect 3299 43 3333 59
rect 4957 119 4991 135
rect 4957 43 4991 59
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect -4991 -121 -4957 -105
rect -4991 -197 -4957 -181
rect -3333 -121 -3299 -105
rect -3333 -197 -3299 -181
rect -1675 -121 -1641 -105
rect -1675 -197 -1641 -181
rect -17 -121 17 -105
rect -17 -197 17 -181
rect 1641 -121 1675 -105
rect 1641 -197 1675 -181
rect 3299 -121 3333 -105
rect 3299 -197 3333 -181
rect 4957 -121 4991 -105
rect 4957 -197 4991 -181
rect -4945 -311 -4929 -277
rect -3361 -311 -3345 -277
rect -3287 -311 -3271 -277
rect -1703 -311 -1687 -277
rect -1629 -311 -1613 -277
rect -45 -311 -29 -277
rect 29 -311 45 -277
rect 1613 -311 1629 -277
rect 1687 -311 1703 -277
rect 3271 -311 3287 -277
rect 3345 -311 3361 -277
rect 4929 -311 4945 -277
rect -4991 -361 -4957 -345
rect -4991 -437 -4957 -421
rect -3333 -361 -3299 -345
rect -3333 -437 -3299 -421
rect -1675 -361 -1641 -345
rect -1675 -437 -1641 -421
rect -17 -361 17 -345
rect -17 -437 17 -421
rect 1641 -361 1675 -345
rect 1641 -437 1675 -421
rect 3299 -361 3333 -345
rect 3299 -437 3333 -421
rect 4957 -361 4991 -345
rect 4957 -437 4991 -421
rect -4945 -551 -4929 -517
rect -3361 -551 -3345 -517
rect -3287 -551 -3271 -517
rect -1703 -551 -1687 -517
rect -1629 -551 -1613 -517
rect -45 -551 -29 -517
rect 29 -551 45 -517
rect 1613 -551 1629 -517
rect 1687 -551 1703 -517
rect 3271 -551 3287 -517
rect 3345 -551 3361 -517
rect 4929 -551 4945 -517
rect -4991 -601 -4957 -585
rect -4991 -677 -4957 -661
rect -3333 -601 -3299 -585
rect -3333 -677 -3299 -661
rect -1675 -601 -1641 -585
rect -1675 -677 -1641 -661
rect -17 -601 17 -585
rect -17 -677 17 -661
rect 1641 -601 1675 -585
rect 1641 -677 1675 -661
rect 3299 -601 3333 -585
rect 3299 -677 3333 -661
rect 4957 -601 4991 -585
rect 4957 -677 4991 -661
rect -4945 -791 -4929 -757
rect -3361 -791 -3345 -757
rect -3287 -791 -3271 -757
rect -1703 -791 -1687 -757
rect -1629 -791 -1613 -757
rect -45 -791 -29 -757
rect 29 -791 45 -757
rect 1613 -791 1629 -757
rect 1687 -791 1703 -757
rect 3271 -791 3287 -757
rect 3345 -791 3361 -757
rect 4929 -791 4945 -757
rect -4991 -841 -4957 -825
rect -4991 -917 -4957 -901
rect -3333 -841 -3299 -825
rect -3333 -917 -3299 -901
rect -1675 -841 -1641 -825
rect -1675 -917 -1641 -901
rect -17 -841 17 -825
rect -17 -917 17 -901
rect 1641 -841 1675 -825
rect 1641 -917 1675 -901
rect 3299 -841 3333 -825
rect 3299 -917 3333 -901
rect 4957 -841 4991 -825
rect 4957 -917 4991 -901
rect -5125 -1027 -5091 -965
rect 5091 -1027 5125 -965
rect -5125 -1061 -5029 -1027
rect 5029 -1061 5125 -1027
<< viali >>
rect -4929 889 -3361 923
rect -3271 889 -1703 923
rect -1613 889 -45 923
rect 45 889 1613 923
rect 1703 889 3271 923
rect 3361 889 4929 923
rect -4991 779 -4957 839
rect -3333 779 -3299 839
rect -1675 779 -1641 839
rect -17 779 17 839
rect 1641 779 1675 839
rect 3299 779 3333 839
rect 4957 779 4991 839
rect -4929 649 -3361 683
rect -3271 649 -1703 683
rect -1613 649 -45 683
rect 45 649 1613 683
rect 1703 649 3271 683
rect 3361 649 4929 683
rect -4991 539 -4957 599
rect -3333 539 -3299 599
rect -1675 539 -1641 599
rect -17 539 17 599
rect 1641 539 1675 599
rect 3299 539 3333 599
rect 4957 539 4991 599
rect -4929 409 -3361 443
rect -3271 409 -1703 443
rect -1613 409 -45 443
rect 45 409 1613 443
rect 1703 409 3271 443
rect 3361 409 4929 443
rect -4991 299 -4957 359
rect -3333 299 -3299 359
rect -1675 299 -1641 359
rect -17 299 17 359
rect 1641 299 1675 359
rect 3299 299 3333 359
rect 4957 299 4991 359
rect -4929 169 -3361 203
rect -3271 169 -1703 203
rect -1613 169 -45 203
rect 45 169 1613 203
rect 1703 169 3271 203
rect 3361 169 4929 203
rect -4991 59 -4957 119
rect -3333 59 -3299 119
rect -1675 59 -1641 119
rect -17 59 17 119
rect 1641 59 1675 119
rect 3299 59 3333 119
rect 4957 59 4991 119
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect -4991 -181 -4957 -121
rect -3333 -181 -3299 -121
rect -1675 -181 -1641 -121
rect -17 -181 17 -121
rect 1641 -181 1675 -121
rect 3299 -181 3333 -121
rect 4957 -181 4991 -121
rect -4929 -311 -3361 -277
rect -3271 -311 -1703 -277
rect -1613 -311 -45 -277
rect 45 -311 1613 -277
rect 1703 -311 3271 -277
rect 3361 -311 4929 -277
rect -4991 -421 -4957 -361
rect -3333 -421 -3299 -361
rect -1675 -421 -1641 -361
rect -17 -421 17 -361
rect 1641 -421 1675 -361
rect 3299 -421 3333 -361
rect 4957 -421 4991 -361
rect -4929 -551 -3361 -517
rect -3271 -551 -1703 -517
rect -1613 -551 -45 -517
rect 45 -551 1613 -517
rect 1703 -551 3271 -517
rect 3361 -551 4929 -517
rect -4991 -661 -4957 -601
rect -3333 -661 -3299 -601
rect -1675 -661 -1641 -601
rect -17 -661 17 -601
rect 1641 -661 1675 -601
rect 3299 -661 3333 -601
rect 4957 -661 4991 -601
rect -4929 -791 -3361 -757
rect -3271 -791 -1703 -757
rect -1613 -791 -45 -757
rect 45 -791 1613 -757
rect 1703 -791 3271 -757
rect 3361 -791 4929 -757
rect -4991 -901 -4957 -841
rect -3333 -901 -3299 -841
rect -1675 -901 -1641 -841
rect -17 -901 17 -841
rect 1641 -901 1675 -841
rect 3299 -901 3333 -841
rect 4957 -901 4991 -841
<< metal1 >>
rect -4997 923 -3349 929
rect -4997 889 -4929 923
rect -3361 889 -3349 923
rect -4997 883 -3349 889
rect -3283 923 -1691 929
rect -3283 889 -3271 923
rect -1703 889 -1691 923
rect -3283 883 -1691 889
rect -1625 923 -33 929
rect -1625 889 -1613 923
rect -45 889 -33 923
rect -1625 883 -33 889
rect 33 923 1625 929
rect 33 889 45 923
rect 1613 889 1625 923
rect 33 883 1625 889
rect 1691 923 3283 929
rect 1691 889 1703 923
rect 3271 889 3283 923
rect 1691 883 3283 889
rect 3349 923 4997 929
rect 3349 889 3361 923
rect 4929 889 4997 923
rect 3349 883 4997 889
rect -4997 839 -4951 883
rect -4997 779 -4991 839
rect -4957 779 -4951 839
rect -4997 767 -4951 779
rect -3339 839 -3293 851
rect -3339 779 -3333 839
rect -3299 779 -3293 839
rect -3339 767 -3293 779
rect -1681 839 -1635 851
rect -1681 779 -1675 839
rect -1641 779 -1635 839
rect -1681 767 -1635 779
rect -23 839 23 851
rect -23 779 -17 839
rect 17 779 23 839
rect -23 767 23 779
rect 1635 839 1681 851
rect 1635 779 1641 839
rect 1675 779 1681 839
rect 1635 767 1681 779
rect 3293 839 3339 851
rect 3293 779 3299 839
rect 3333 779 3339 839
rect 3293 767 3339 779
rect 4951 839 4997 883
rect 4951 779 4957 839
rect 4991 779 4997 839
rect 4951 767 4997 779
rect -4997 683 -3349 689
rect -4997 649 -4929 683
rect -3361 649 -3349 683
rect -4997 643 -3349 649
rect -3283 683 -1691 689
rect -3283 649 -3271 683
rect -1703 649 -1691 683
rect -3283 643 -1691 649
rect -1625 683 -33 689
rect -1625 649 -1613 683
rect -45 649 -33 683
rect -1625 643 -33 649
rect 33 683 1625 689
rect 33 649 45 683
rect 1613 649 1625 683
rect 33 643 1625 649
rect 1691 683 3283 689
rect 1691 649 1703 683
rect 3271 649 3283 683
rect 1691 643 3283 649
rect 3349 683 4997 689
rect 3349 649 3361 683
rect 4929 649 4997 683
rect 3349 643 4997 649
rect -4997 599 -4951 643
rect -4997 539 -4991 599
rect -4957 539 -4951 599
rect -4997 527 -4951 539
rect -3339 599 -3293 611
rect -3339 539 -3333 599
rect -3299 539 -3293 599
rect -3339 527 -3293 539
rect -1681 599 -1635 611
rect -1681 539 -1675 599
rect -1641 539 -1635 599
rect -1681 527 -1635 539
rect -23 599 23 611
rect -23 539 -17 599
rect 17 539 23 599
rect -23 527 23 539
rect 1635 599 1681 611
rect 1635 539 1641 599
rect 1675 539 1681 599
rect 1635 527 1681 539
rect 3293 599 3339 611
rect 3293 539 3299 599
rect 3333 539 3339 599
rect 3293 527 3339 539
rect 4951 599 4997 643
rect 4951 539 4957 599
rect 4991 539 4997 599
rect 4951 527 4997 539
rect -4997 443 -3349 449
rect -4997 409 -4929 443
rect -3361 409 -3349 443
rect -4997 403 -3349 409
rect -3283 443 -1691 449
rect -3283 409 -3271 443
rect -1703 409 -1691 443
rect -3283 403 -1691 409
rect -1625 443 -33 449
rect -1625 409 -1613 443
rect -45 409 -33 443
rect -1625 403 -33 409
rect 33 443 1625 449
rect 33 409 45 443
rect 1613 409 1625 443
rect 33 403 1625 409
rect 1691 443 3283 449
rect 1691 409 1703 443
rect 3271 409 3283 443
rect 1691 403 3283 409
rect 3349 443 4997 449
rect 3349 409 3361 443
rect 4929 409 4997 443
rect 3349 403 4997 409
rect -4997 359 -4951 403
rect -4997 299 -4991 359
rect -4957 299 -4951 359
rect -4997 287 -4951 299
rect -3339 359 -3293 371
rect -3339 299 -3333 359
rect -3299 299 -3293 359
rect -3339 287 -3293 299
rect -1681 359 -1635 371
rect -1681 299 -1675 359
rect -1641 299 -1635 359
rect -1681 287 -1635 299
rect -23 359 23 371
rect -23 299 -17 359
rect 17 299 23 359
rect -23 287 23 299
rect 1635 359 1681 371
rect 1635 299 1641 359
rect 1675 299 1681 359
rect 1635 287 1681 299
rect 3293 359 3339 371
rect 3293 299 3299 359
rect 3333 299 3339 359
rect 3293 287 3339 299
rect 4951 359 4997 403
rect 4951 299 4957 359
rect 4991 299 4997 359
rect 4951 287 4997 299
rect -4997 203 -3349 209
rect -4997 169 -4929 203
rect -3361 169 -3349 203
rect -4997 163 -3349 169
rect -3283 203 -1691 209
rect -3283 169 -3271 203
rect -1703 169 -1691 203
rect -3283 163 -1691 169
rect -1625 203 -33 209
rect -1625 169 -1613 203
rect -45 169 -33 203
rect -1625 163 -33 169
rect 33 203 1625 209
rect 33 169 45 203
rect 1613 169 1625 203
rect 33 163 1625 169
rect 1691 203 3283 209
rect 1691 169 1703 203
rect 3271 169 3283 203
rect 1691 163 3283 169
rect 3349 203 4997 209
rect 3349 169 3361 203
rect 4929 169 4997 203
rect 3349 163 4997 169
rect -4997 119 -4951 163
rect -4997 59 -4991 119
rect -4957 59 -4951 119
rect -4997 47 -4951 59
rect -3339 119 -3293 131
rect -3339 59 -3333 119
rect -3299 59 -3293 119
rect -3339 47 -3293 59
rect -1681 119 -1635 131
rect -1681 59 -1675 119
rect -1641 59 -1635 119
rect -1681 47 -1635 59
rect -23 119 23 131
rect -23 59 -17 119
rect 17 59 23 119
rect -23 47 23 59
rect 1635 119 1681 131
rect 1635 59 1641 119
rect 1675 59 1681 119
rect 1635 47 1681 59
rect 3293 119 3339 131
rect 3293 59 3299 119
rect 3333 59 3339 119
rect 3293 47 3339 59
rect 4951 119 4997 163
rect 4951 59 4957 119
rect 4991 59 4997 119
rect 4951 47 4997 59
rect -4997 -37 -3349 -31
rect -4997 -71 -4929 -37
rect -3361 -71 -3349 -37
rect -4997 -77 -3349 -71
rect -3283 -37 -1691 -31
rect -3283 -71 -3271 -37
rect -1703 -71 -1691 -37
rect -3283 -77 -1691 -71
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect 1691 -37 3283 -31
rect 1691 -71 1703 -37
rect 3271 -71 3283 -37
rect 1691 -77 3283 -71
rect 3349 -37 4997 -31
rect 3349 -71 3361 -37
rect 4929 -71 4997 -37
rect 3349 -77 4997 -71
rect -4997 -121 -4951 -77
rect -4997 -181 -4991 -121
rect -4957 -181 -4951 -121
rect -4997 -193 -4951 -181
rect -3339 -121 -3293 -109
rect -3339 -181 -3333 -121
rect -3299 -181 -3293 -121
rect -3339 -193 -3293 -181
rect -1681 -121 -1635 -109
rect -1681 -181 -1675 -121
rect -1641 -181 -1635 -121
rect -1681 -193 -1635 -181
rect -23 -121 23 -109
rect -23 -181 -17 -121
rect 17 -181 23 -121
rect -23 -193 23 -181
rect 1635 -121 1681 -109
rect 1635 -181 1641 -121
rect 1675 -181 1681 -121
rect 1635 -193 1681 -181
rect 3293 -121 3339 -109
rect 3293 -181 3299 -121
rect 3333 -181 3339 -121
rect 3293 -193 3339 -181
rect 4951 -121 4997 -77
rect 4951 -181 4957 -121
rect 4991 -181 4997 -121
rect 4951 -193 4997 -181
rect -4997 -277 -3349 -271
rect -4997 -311 -4929 -277
rect -3361 -311 -3349 -277
rect -4997 -317 -3349 -311
rect -3283 -277 -1691 -271
rect -3283 -311 -3271 -277
rect -1703 -311 -1691 -277
rect -3283 -317 -1691 -311
rect -1625 -277 -33 -271
rect -1625 -311 -1613 -277
rect -45 -311 -33 -277
rect -1625 -317 -33 -311
rect 33 -277 1625 -271
rect 33 -311 45 -277
rect 1613 -311 1625 -277
rect 33 -317 1625 -311
rect 1691 -277 3283 -271
rect 1691 -311 1703 -277
rect 3271 -311 3283 -277
rect 1691 -317 3283 -311
rect 3349 -277 4997 -271
rect 3349 -311 3361 -277
rect 4929 -311 4997 -277
rect 3349 -317 4997 -311
rect -4997 -361 -4951 -317
rect -4997 -421 -4991 -361
rect -4957 -421 -4951 -361
rect -4997 -433 -4951 -421
rect -3339 -361 -3293 -349
rect -3339 -421 -3333 -361
rect -3299 -421 -3293 -361
rect -3339 -433 -3293 -421
rect -1681 -361 -1635 -349
rect -1681 -421 -1675 -361
rect -1641 -421 -1635 -361
rect -1681 -433 -1635 -421
rect -23 -361 23 -349
rect -23 -421 -17 -361
rect 17 -421 23 -361
rect -23 -433 23 -421
rect 1635 -361 1681 -349
rect 1635 -421 1641 -361
rect 1675 -421 1681 -361
rect 1635 -433 1681 -421
rect 3293 -361 3339 -349
rect 3293 -421 3299 -361
rect 3333 -421 3339 -361
rect 3293 -433 3339 -421
rect 4951 -361 4997 -317
rect 4951 -421 4957 -361
rect 4991 -421 4997 -361
rect 4951 -433 4997 -421
rect -4997 -517 -3349 -511
rect -4997 -551 -4929 -517
rect -3361 -551 -3349 -517
rect -4997 -557 -3349 -551
rect -3283 -517 -1691 -511
rect -3283 -551 -3271 -517
rect -1703 -551 -1691 -517
rect -3283 -557 -1691 -551
rect -1625 -517 -33 -511
rect -1625 -551 -1613 -517
rect -45 -551 -33 -517
rect -1625 -557 -33 -551
rect 33 -517 1625 -511
rect 33 -551 45 -517
rect 1613 -551 1625 -517
rect 33 -557 1625 -551
rect 1691 -517 3283 -511
rect 1691 -551 1703 -517
rect 3271 -551 3283 -517
rect 1691 -557 3283 -551
rect 3349 -517 4997 -511
rect 3349 -551 3361 -517
rect 4929 -551 4997 -517
rect 3349 -557 4997 -551
rect -4997 -601 -4951 -557
rect -4997 -661 -4991 -601
rect -4957 -661 -4951 -601
rect -4997 -673 -4951 -661
rect -3339 -601 -3293 -589
rect -3339 -661 -3333 -601
rect -3299 -661 -3293 -601
rect -3339 -673 -3293 -661
rect -1681 -601 -1635 -589
rect -1681 -661 -1675 -601
rect -1641 -661 -1635 -601
rect -1681 -673 -1635 -661
rect -23 -601 23 -589
rect -23 -661 -17 -601
rect 17 -661 23 -601
rect -23 -673 23 -661
rect 1635 -601 1681 -589
rect 1635 -661 1641 -601
rect 1675 -661 1681 -601
rect 1635 -673 1681 -661
rect 3293 -601 3339 -589
rect 3293 -661 3299 -601
rect 3333 -661 3339 -601
rect 3293 -673 3339 -661
rect 4951 -601 4997 -557
rect 4951 -661 4957 -601
rect 4991 -661 4997 -601
rect 4951 -673 4997 -661
rect -4997 -757 -3349 -751
rect -4997 -791 -4929 -757
rect -3361 -791 -3349 -757
rect -4997 -797 -3349 -791
rect -3283 -757 -1691 -751
rect -3283 -791 -3271 -757
rect -1703 -791 -1691 -757
rect -3283 -797 -1691 -791
rect -1625 -757 -33 -751
rect -1625 -791 -1613 -757
rect -45 -791 -33 -757
rect -1625 -797 -33 -791
rect 33 -757 1625 -751
rect 33 -791 45 -757
rect 1613 -791 1625 -757
rect 33 -797 1625 -791
rect 1691 -757 3283 -751
rect 1691 -791 1703 -757
rect 3271 -791 3283 -757
rect 1691 -797 3283 -791
rect 3349 -757 4997 -751
rect 3349 -791 3361 -757
rect 4929 -791 4997 -757
rect 3349 -797 4997 -791
rect -4997 -841 -4951 -797
rect -4997 -901 -4991 -841
rect -4957 -901 -4951 -841
rect -4997 -913 -4951 -901
rect -3339 -841 -3293 -829
rect -3339 -901 -3333 -841
rect -3299 -901 -3293 -841
rect -3339 -913 -3293 -901
rect -1681 -841 -1635 -829
rect -1681 -901 -1675 -841
rect -1641 -901 -1635 -841
rect -1681 -913 -1635 -901
rect -23 -841 23 -829
rect -23 -901 -17 -841
rect 17 -901 23 -841
rect -23 -913 23 -901
rect 1635 -841 1681 -829
rect 1635 -901 1641 -841
rect 1675 -901 1681 -841
rect 1635 -913 1681 -901
rect 3293 -841 3339 -829
rect 3293 -901 3299 -841
rect 3333 -901 3339 -841
rect 3293 -913 3339 -901
rect 4951 -841 4997 -797
rect 4951 -901 4957 -841
rect 4991 -901 4997 -841
rect 4951 -913 4997 -901
<< metal2 >>
rect -5000 -839 -4948 777
rect -3342 -839 -3290 777
rect -1684 -839 -1632 777
rect -26 -839 26 777
rect 1632 -839 1684 777
rect 3290 -839 3342 777
rect 4948 -839 5000 777
<< properties >>
string FIXED_BBOX -5108 -1044 5108 1044
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 8 m 8 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
* NGSPICE file created from brownout_dig.ext - technology: sky130A
* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt brownout_dig a_VGND a_VPWR a_brout_filt a_ena a_force_rc_osc a_force_short_oneshot a_osc_ck a_osc_ck_256 a_osc_ena a_otrip_0_ a_otrip_1_ a_otrip_2_ a_otrip_decoded_0_ a_otrip_decoded_1_ a_otrip_decoded_2_ a_otrip_decoded_3_ a_otrip_decoded_4_ a_otrip_decoded_5_ a_otrip_decoded_6_ a_otrip_decoded_7_ a_out_unbuf a_timed_out a_vtrip_0_ a_vtrip_1_ a_vtrip_2_ a_vtrip_decoded_0_ a_vtrip_decoded_1_ a_vtrip_decoded_2_ a_vtrip_decoded_3_ a_vtrip_decoded_4_ a_vtrip_decoded_5_ a_vtrip_decoded_6_ a_vtrip_decoded_7_
A_131_ [cnt\_10\_ net31] _049_ d_lut_sky130_fd_sc_hd__or2_1
A_114_ [_033_ _038_ net32] _010_ d_lut_sky130_fd_sc_hd__a21oi_1
Aoutput20 [net20] otrip_decoded_7_ d_lut_sky130_fd_sc_hd__clkbuf_4
A_130_ [cnt\_9\_ cnt\_8\_ _067_ net4] _048_ d_lut_sky130_fd_sc_hd__a31o_1
Aclkbuf_2_3__f_osc_ck [clknet_0_osc_ck] clknet_2_3__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_113_ [_063_ _037_] _038_ d_lut_sky130_fd_sc_hd__nand2b_1
Aoutput21 [net21] out_unbuf d_lut_sky130_fd_sc_hd__buf_2
A_189_ _005_ clknet_2_2__leaf_osc_ck NULL ~net37 cnt_ck_256\_5\_ NULL ddflop
A_112_ [cnt\_1\_ cnt\_0\_ cnt\_2\_ cnt\_3\_] _037_ d_lut_sky130_fd_sc_hd__a31o_1
Ahold10 [cnt_ck_256\_1\_] net46 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput22 [net22] timed_out d_lut_sky130_fd_sc_hd__buf_2
Aoutput11 [net11] osc_ck_256 d_lut_sky130_fd_sc_hd__buf_2
A_188_ _004_ clknet_2_2__leaf_osc_ck NULL ~net37 cnt_ck_256\_4\_ NULL ddflop
A_111_ [_033_ _036_ net43] _009_ d_lut_sky130_fd_sc_hd__a21oi_1
Ahold11 [_001_] net47 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput12 [net12] osc_ena d_lut_sky130_fd_sc_hd__buf_2
Aoutput23 [net23] vtrip_decoded_0_ d_lut_sky130_fd_sc_hd__buf_2
A_187_ _003_ clknet_2_2__leaf_osc_ck NULL ~net37 cnt_ck_256\_3\_ NULL ddflop
A_110_ [cnt\_2\_ _062_] _036_ d_lut_sky130_fd_sc_hd__xor2_1
Ahold12 [cnt_ck_256\_0\_] net48 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput24 [net24] vtrip_decoded_1_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput13 [net13] otrip_decoded_0_ d_lut_sky130_fd_sc_hd__buf_2
A_186_ _002_ clknet_2_3__leaf_osc_ck NULL ~net37 cnt_ck_256\_2\_ NULL ddflop
A_169_ _008_ clknet_2_3__leaf_osc_ck ~net34 NULL cnt\_1\_ NULL ddflop
Ahold13 [cnt_ck_256\_5\_] net49 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput25 [net25] vtrip_decoded_2_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput14 [net14] otrip_decoded_1_ d_lut_sky130_fd_sc_hd__buf_2
A_185_ net47 clknet_2_3__leaf_osc_ck NULL ~net37 cnt_ck_256\_1\_ NULL ddflop
A_168_ _007_ clknet_2_3__leaf_osc_ck ~net34 NULL cnt\_0\_ NULL ddflop
A_099_ [cnt_ck_256\_5\_ cnt_ck_256\_4\_ _027_] _029_ d_lut_sky130_fd_sc_hd__and3_1
Ahold14 [_030_] net50 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput26 [net26] vtrip_decoded_3_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput15 [net15] otrip_decoded_2_ d_lut_sky130_fd_sc_hd__buf_2
A_184_ _000_ clknet_2_3__leaf_osc_ck NULL ~net37 cnt_ck_256\_0\_ NULL ddflop
A_098_ [net51 _027_] _004_ d_lut_sky130_fd_sc_hd__xor2_1
A_167_ [net7 net6 net5] net14 d_lut_sky130_fd_sc_hd__nor3b_1
Ahold15 [cnt_ck_256\_4\_] net51 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput16 [net16] otrip_decoded_3_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput27 [net27] vtrip_decoded_4_ d_lut_sky130_fd_sc_hd__buf_2
A_183_ _022_ clknet_2_0__leaf_osc_ck ~net33 NULL cnt\_15\_ NULL ddflop
A_097_ [_027_ _028_] _003_ d_lut_sky130_fd_sc_hd__nor2_1
A_166_ [net7 net5 net6] net13 d_lut_sky130_fd_sc_hd__nor3_1
Ahold16 [cnt_ck_256\_2\_] net52 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_149_ [net45 _031_] _023_ d_lut_sky130_fd_sc_hd__xnor2_1
Aoutput17 [net17] otrip_decoded_4_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput28 [net28] vtrip_decoded_5_ d_lut_sky130_fd_sc_hd__buf_2
A_182_ _021_ clknet_2_0__leaf_osc_ck ~net33 NULL cnt\_14\_ NULL ddflop
A_165_ [_073_] net21 d_lut_sky130_fd_sc_hd__inv_2
A_096_ [net53 _025_] _028_ d_lut_sky130_fd_sc_hd__nor2_1
Ahold17 [cnt_ck_256\_3\_] net53 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_148_ [_061_ _059_ _060_ _024_] _022_ d_lut_sky130_fd_sc_hd__a31o_1
A_079_ [net7 net5 net6] net20 d_lut_sky130_fd_sc_hd__and3_1
Aoutput29 [net29] vtrip_decoded_6_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput18 [net18] otrip_decoded_5_ d_lut_sky130_fd_sc_hd__buf_2
Aclkbuf_2_2__f_osc_ck [clknet_0_osc_ck] clknet_2_2__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
Afanout31 [_048_] net31 d_lut_sky130_fd_sc_hd__clkbuf_2
A_181_ _020_ clknet_2_1__leaf_osc_ck ~net33 NULL cnt\_13\_ NULL ddflop
A_164_ [_061_ net22] _073_ d_lut_sky130_fd_sc_hd__nand2_1
A_095_ [cnt_ck_256\_3\_ _025_] _027_ d_lut_sky130_fd_sc_hd__and2_1
A_147_ [cnt\_15\_ _071_ net31] _060_ d_lut_sky130_fd_sc_hd__nand3_1
A_078_ [net5 net6 net7] net19 d_lut_sky130_fd_sc_hd__and3b_1
Aoutput19 [net19] otrip_decoded_6_ d_lut_sky130_fd_sc_hd__buf_2
A_180_ _019_ clknet_2_3__leaf_osc_ck ~net33 NULL cnt\_12\_ NULL ddflop
Afanout32 [brout_filt_retimed] net32 d_lut_sky130_fd_sc_hd__buf_2
A_163_ [cnt\_9\_ cnt\_8\_ _067_ _072_] net22 d_lut_sky130_fd_sc_hd__and4_1
A_094_ [_025_ _026_] _002_ d_lut_sky130_fd_sc_hd__nor2_1
A_077_ [net6 net5 net7] net18 d_lut_sky130_fd_sc_hd__and3b_1
A_146_ [_071_ net31 cnt\_15\_] _059_ d_lut_sky130_fd_sc_hd__a21o_1
A_129_ [_033_ _047_ net32] _016_ d_lut_sky130_fd_sc_hd__a21oi_1
Afanout33 [net42] net33 d_lut_sky130_fd_sc_hd__clkbuf_4
A_162_ [cnt\_14\_ cnt\_15\_ _070_] _072_ d_lut_sky130_fd_sc_hd__and3_1
A_093_ [cnt_ck_256\_0\_ net46 net52] _026_ d_lut_sky130_fd_sc_hd__a21oi_1
Ainput1 [brout_filt] net1 d_lut_sky130_fd_sc_hd__clkbuf_1
A_145_ [_061_ _057_ _058_ _024_] _021_ d_lut_sky130_fd_sc_hd__a31o_1
A_076_ [net5 net6 net7] net17 d_lut_sky130_fd_sc_hd__nor3b_1
A_128_ [_068_ _046_] _047_ d_lut_sky130_fd_sc_hd__or2_1
Afanout34 [net42] net34 d_lut_sky130_fd_sc_hd__clkbuf_2
A_161_ [cnt\_14\_ _070_] _071_ d_lut_sky130_fd_sc_hd__and2_1
A_092_ [cnt_ck_256\_0\_ cnt_ck_256\_1\_ cnt_ck_256\_2\_] _025_ d_lut_sky130_fd_sc_hd__and3_1
Ainput2 [ena] net2 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_075_ [net7 net5 net6] net16 d_lut_sky130_fd_sc_hd__and3b_1
A_144_ [_071_ net31] _058_ d_lut_sky130_fd_sc_hd__nand2_1
A_197__360 net36 done
A_197__361 _197__36/LO dzero
A_127_ [cnt\_8\_ _067_ cnt\_9\_] _046_ d_lut_sky130_fd_sc_hd__a21oi_1
A_160_ [cnt\_11\_ cnt\_10\_ cnt\_13\_ cnt\_12\_] _070_ d_lut_sky130_fd_sc_hd__and4_1
A_091_ [cnt_ck_256\_0\_ net46] _001_ d_lut_sky130_fd_sc_hd__xor2_1
Ainput3 [force_rc_osc] net3 d_lut_sky130_fd_sc_hd__clkbuf_1
A_143_ [_070_ net31 cnt\_14\_] _057_ d_lut_sky130_fd_sc_hd__a21o_1
A_074_ [net7 net5 net6] net15 d_lut_sky130_fd_sc_hd__nor3b_1
A_126_ [_033_ _045_ net32] _015_ d_lut_sky130_fd_sc_hd__a21oi_1
A_109_ [_033_ _035_ net43] _008_ d_lut_sky130_fd_sc_hd__a21oi_1
A_090_ [net2 _073_ brout_filt_ena_rsb net3] net12 d_lut_sky130_fd_sc_hd__a211o_1
Ainput4 [force_short_oneshot] net4 d_lut_sky130_fd_sc_hd__buf_1
A_142_ [_055_ _056_ _024_] _020_ d_lut_sky130_fd_sc_hd__a21o_1
A_125_ [cnt\_8\_ _067_] _045_ d_lut_sky130_fd_sc_hd__xnor2_1
A_108_ [_062_ _034_] _035_ d_lut_sky130_fd_sc_hd__nand2_1
Ainput5 [otrip_0_] net5 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_141_ [_070_ _048_ net32] _056_ d_lut_sky130_fd_sc_hd__a21oi_1
A_124_ [_033_ _044_ net32] _014_ d_lut_sky130_fd_sc_hd__a21oi_1
A_107_ [cnt\_1\_ cnt\_0\_] _034_ d_lut_sky130_fd_sc_hd__or2_1
Ainput6 [otrip_1_] net6 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_140_ [_069_ _048_ cnt\_13\_] _055_ d_lut_sky130_fd_sc_hd__a21o_1
A_123_ [cnt\_7\_ _066_] _044_ d_lut_sky130_fd_sc_hd__xnor2_1
A_106_ [net44 _033_ net43] _007_ d_lut_sky130_fd_sc_hd__a21oi_1
Ainput7 [otrip_2_] net7 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_122_ [_033_ _043_ net32] _013_ d_lut_sky130_fd_sc_hd__a21oi_1
Ainput10 [vtrip_2_] net10 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
Aclkbuf_2_1__f_osc_ck [clknet_0_osc_ck] clknet_2_1__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_105_ [net4 net22] _033_ d_lut_sky130_fd_sc_hd__nor2_2
Ainput8 [vtrip_0_] net8 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_198_ net39 clknet_2_2__leaf_osc_ck NULL ~brout_filt_ena_rsb brout_filt_retime_rsb NULL ddflop
A_121_ [_066_ _042_] _043_ d_lut_sky130_fd_sc_hd__nand2b_1
A_104_ [_031_ _032_] _006_ d_lut_sky130_fd_sc_hd__and2_1
Ainput9 [vtrip_1_] net9 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_197_ net36 clknet_2_0__leaf_osc_ck NULL ~brout_filt_ena_rsb brout_filt_retime_rsb_stg1 NULL ddflop
A_120_ [cnt\_5\_ cnt\_4\_ _063_ cnt\_6\_] _042_ d_lut_sky130_fd_sc_hd__a31o_1
A_103_ [cnt_ck_256\_6\_ _029_] _032_ d_lut_sky130_fd_sc_hd__or2_1
Ahold1 [brout_filt_retime_rsb] net37 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_196_ net38 clknet_2_2__leaf_osc_ck NULL ~net37 brout_filt_retimed NULL ddflop
A_179_ _018_ clknet_2_2__leaf_osc_ck ~net33 NULL cnt\_11\_ NULL ddflop
Aclkbuf_0_osc_ck [osc_ck] clknet_0_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_102_ [cnt_ck_256\_6\_ _029_] _031_ d_lut_sky130_fd_sc_hd__nand2_1
Ahold2 [brout_filt_retimed_stg1] net38 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_195_ net1 clknet_2_0__leaf_osc_ck NULL ~net37 brout_filt_retimed_stg1 NULL ddflop
A_178_ _017_ clknet_2_2__leaf_osc_ck ~net33 NULL cnt\_10\_ NULL ddflop
A_101_ [_029_ net50] _005_ d_lut_sky130_fd_sc_hd__nor2_1
Ahold3 [brout_filt_retime_rsb_stg1] net39 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_194_ net41 clknet_2_0__leaf_osc_ck NULL ~net2 cnt_rsb NULL ddflop
A_177_ _016_ clknet_2_1__leaf_osc_ck ~net33 NULL cnt\_9\_ NULL ddflop
A_100_ [cnt_ck_256\_4\_ _027_ net49] _030_ d_lut_sky130_fd_sc_hd__a21oi_1
Ahold4 [cnt_rsb_stg1] net40 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_193_ net40 clknet_2_0__leaf_osc_ck NULL ~net2 cnt_rsb_stg2 NULL ddflop
A_176_ _015_ clknet_2_1__leaf_osc_ck ~net33 NULL cnt\_8\_ NULL ddflop
A_159_ [cnt\_11\_ cnt\_10\_ cnt\_12\_] _069_ d_lut_sky130_fd_sc_hd__and3_1
Ahold5 [cnt_rsb_stg2] net41 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_192_ net35 clknet_2_0__leaf_osc_ck NULL ~net2 cnt_rsb_stg1 NULL ddflop
A_175_ _014_ clknet_2_1__leaf_osc_ck ~net33 NULL cnt\_7\_ NULL ddflop
A_158_ [cnt\_9\_ cnt\_8\_ _067_] _068_ d_lut_sky130_fd_sc_hd__and3_1
A_089_ [net1 net2] brout_filt_ena_rsb d_lut_sky130_fd_sc_hd__and2_1
Ahold6 [cnt_rsb] net42 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_191_ _023_ clknet_2_2__leaf_osc_ck NULL ~net37 net11 NULL ddflop
A_174_ _013_ clknet_2_1__leaf_osc_ck ~net33 NULL cnt\_6\_ NULL ddflop
A_157_ [cnt\_4\_ cnt\_7\_ _063_ _065_] _067_ d_lut_sky130_fd_sc_hd__and4_1
A_088_ [_061_ cnt\_15\_ _068_ _071_] _024_ d_lut_sky130_fd_sc_hd__and4_2
Ahold7 [brout_filt_retimed] net43 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aclkbuf_2_0__f_osc_ck [clknet_0_osc_ck] clknet_2_0__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_190_ _006_ clknet_2_2__leaf_osc_ck NULL ~net37 cnt_ck_256\_6\_ NULL ddflop
A_173_ _012_ clknet_2_1__leaf_osc_ck ~net34 NULL cnt\_5\_ NULL ddflop
A_156_ [cnt\_4\_ _063_ _065_] _066_ d_lut_sky130_fd_sc_hd__and3_1
A_087_ [net10 net9 net8] net30 d_lut_sky130_fd_sc_hd__and3_1
Ahold8 [cnt\_0\_] net44 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_139_ [_053_ _054_ _024_] _019_ d_lut_sky130_fd_sc_hd__a21o_1
A_172_ _011_ clknet_2_1__leaf_osc_ck ~net34 NULL cnt\_4\_ NULL ddflop
A_086_ [net8 net9 net10] net29 d_lut_sky130_fd_sc_hd__and3b_1
A_155_ [cnt\_5\_ cnt\_6\_] _065_ d_lut_sky130_fd_sc_hd__and2_1
Ahold9 [net11] net45 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_138_ [_069_ net31 net32] _054_ d_lut_sky130_fd_sc_hd__a21oi_1
A_171_ _010_ clknet_2_3__leaf_osc_ck ~net34 NULL cnt\_3\_ NULL ddflop
A_085_ [net9 net8 net10] net28 d_lut_sky130_fd_sc_hd__and3b_1
A_154_ [cnt\_4\_ _063_] _064_ d_lut_sky130_fd_sc_hd__nand2_1
A_137_ [cnt\_11\_ cnt\_10\_ net31 cnt\_12\_] _053_ d_lut_sky130_fd_sc_hd__a31o_1
A_170_ _009_ clknet_2_3__leaf_osc_ck ~net34 NULL cnt\_2\_ NULL ddflop
A_084_ [net9 net8 net10] net27 d_lut_sky130_fd_sc_hd__nor3b_1
A_153_ [cnt\_1\_ cnt\_0\_ cnt\_3\_ cnt\_2\_] _063_ d_lut_sky130_fd_sc_hd__and4_1
A_136_ [_061_ _051_ _052_ _024_] _018_ d_lut_sky130_fd_sc_hd__a31o_1
A_119_ [_033_ _041_ net32] _012_ d_lut_sky130_fd_sc_hd__a21oi_1
A_192__350 net35 done
A_192__351 _192__35/LO dzero
A_083_ [net10 net9 net8] net26 d_lut_sky130_fd_sc_hd__and3b_1
A_152_ [cnt\_1\_ cnt\_0\_] _062_ d_lut_sky130_fd_sc_hd__nand2_1
A_135_ [cnt\_11\_ cnt\_10\_ net31] _052_ d_lut_sky130_fd_sc_hd__nand3_1
A_118_ [cnt\_5\_ _064_] _041_ d_lut_sky130_fd_sc_hd__xor2_1
A_082_ [net10 net8 net9] net25 d_lut_sky130_fd_sc_hd__nor3b_1
A_151_ [net32] _061_ d_lut_sky130_fd_sc_hd__inv_2
A_134_ [cnt\_10\_ net31 cnt\_11\_] _051_ d_lut_sky130_fd_sc_hd__a21o_1
A_117_ [_033_ _040_ net32] _011_ d_lut_sky130_fd_sc_hd__a21oi_1
A_081_ [net10 net9 net8] net24 d_lut_sky130_fd_sc_hd__nor3b_1
A_150_ [net48] _000_ d_lut_sky130_fd_sc_hd__inv_2
A_133_ [_061_ _049_ _050_ _024_] _017_ d_lut_sky130_fd_sc_hd__a31o_1
A_116_ [_064_ _039_] _040_ d_lut_sky130_fd_sc_hd__nand2_1
A_080_ [net10 net9 net8] net23 d_lut_sky130_fd_sc_hd__nor3_1
A_132_ [cnt\_10\_ net31] _050_ d_lut_sky130_fd_sc_hd__nand2_1
A_115_ [cnt\_4\_ _063_] _039_ d_lut_sky130_fd_sc_hd__or2_1
Aoutput30 [net30] vtrip_decoded_7_ d_lut_sky130_fd_sc_hd__buf_2

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dlatch d_dlatch(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_VGND] [VGND] todig_1v8
AA2D2 [a_VPWR] [VPWR] todig_1v8
AA2D3 [a_brout_filt] [brout_filt] todig_1v8
AA2D4 [a_ena] [ena] todig_1v8
AA2D5 [a_force_rc_osc] [force_rc_osc] todig_1v8
AA2D6 [a_force_short_oneshot] [force_short_oneshot] todig_1v8
AA2D7 [a_osc_ck] [osc_ck] todig_1v8
AD2A1 [osc_ck_256] [a_osc_ck_256] toana_1v8
AD2A2 [osc_ena] [a_osc_ena] toana_1v8
AA2D8 [a_otrip_0_] [otrip_0_] todig_1v8
AA2D9 [a_otrip_1_] [otrip_1_] todig_1v8
AA2D10 [a_otrip_2_] [otrip_2_] todig_1v8
AD2A3 [otrip_decoded_0_] [a_otrip_decoded_0_] toana_1v8
AD2A4 [otrip_decoded_1_] [a_otrip_decoded_1_] toana_1v8
AD2A5 [otrip_decoded_2_] [a_otrip_decoded_2_] toana_1v8
AD2A6 [otrip_decoded_3_] [a_otrip_decoded_3_] toana_1v8
AD2A7 [otrip_decoded_4_] [a_otrip_decoded_4_] toana_1v8
AD2A8 [otrip_decoded_5_] [a_otrip_decoded_5_] toana_1v8
AD2A9 [otrip_decoded_6_] [a_otrip_decoded_6_] toana_1v8
AD2A10 [otrip_decoded_7_] [a_otrip_decoded_7_] toana_1v8
AD2A11 [out_unbuf] [a_out_unbuf] toana_1v8
AD2A12 [timed_out] [a_timed_out] toana_1v8
AA2D11 [a_vtrip_0_] [vtrip_0_] todig_1v8
AA2D12 [a_vtrip_1_] [vtrip_1_] todig_1v8
AA2D13 [a_vtrip_2_] [vtrip_2_] todig_1v8
AD2A13 [vtrip_decoded_0_] [a_vtrip_decoded_0_] toana_1v8
AD2A14 [vtrip_decoded_1_] [a_vtrip_decoded_1_] toana_1v8
AD2A15 [vtrip_decoded_2_] [a_vtrip_decoded_2_] toana_1v8
AD2A16 [vtrip_decoded_3_] [a_vtrip_decoded_3_] toana_1v8
AD2A17 [vtrip_decoded_4_] [a_vtrip_decoded_4_] toana_1v8
AD2A18 [vtrip_decoded_5_] [a_vtrip_decoded_5_] toana_1v8
AD2A19 [vtrip_decoded_6_] [a_vtrip_decoded_6_] toana_1v8
AD2A20 [vtrip_decoded_7_] [a_vtrip_decoded_7_] toana_1v8

.ends


* sky130_ef_sc_hd__decap_12 (no function)
* sky130_fd_sc_hd__or2_1 (A) | (B)
.model d_lut_sky130_fd_sc_hd__or2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0111")
* sky130_fd_sc_hd__decap_8 (no function)
* sky130_fd_sc_hd__a21oi_1 (!A1&!B1) | (!A2&!B1)
.model d_lut_sky130_fd_sc_hd__a21oi_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11100000")
* sky130_fd_sc_hd__fill_1 (no function)
* sky130_fd_sc_hd__tapvpwrvgnd_1 (no function)
* sky130_fd_sc_hd__decap_3 (no function)
* sky130_fd_sc_hd__clkbuf_4 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_4 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__a31o_1 (A1&A2&A3) | (B1)
.model d_lut_sky130_fd_sc_hd__a31o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000111111111")
* sky130_fd_sc_hd__decap_6 (no function)
* sky130_fd_sc_hd__decap_4 (no function)
* sky130_fd_sc_hd__clkbuf_16 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_16 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__nand2b_1 (A_N) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1101")
* sky130_fd_sc_hd__buf_2 (A)
.model d_lut_sky130_fd_sc_hd__buf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__dfrtp_1 IQ
* sky130_fd_sc_hd__fill_2 (no function)
* sky130_fd_sc_hd__dlygate4sd3_1 (A)
.model d_lut_sky130_fd_sc_hd__dlygate4sd3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__xor2_1 (A&!B) | (!A&B)
.model d_lut_sky130_fd_sc_hd__xor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0110")
* sky130_fd_sc_hd__dfstp_1 IQ
* sky130_fd_sc_hd__and3_1 (A&B&C)
.model d_lut_sky130_fd_sc_hd__and3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000001")
* sky130_fd_sc_hd__nor3b_1 (!A&!B&C_N)
.model d_lut_sky130_fd_sc_hd__nor3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00001000")
* sky130_fd_sc_hd__nor2_1 (!A&!B)
.model d_lut_sky130_fd_sc_hd__nor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1000")
* sky130_fd_sc_hd__nor3_1 (!A&!B&!C)
.model d_lut_sky130_fd_sc_hd__nor3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10000000")
* sky130_fd_sc_hd__xnor2_1 (!A&!B) | (A&B)
.model d_lut_sky130_fd_sc_hd__xnor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1001")
* sky130_fd_sc_hd__inv_2 (!A)
.model d_lut_sky130_fd_sc_hd__inv_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10")
* sky130_fd_sc_hd__clkbuf_2 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__nand2_1 (!A) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1110")
* sky130_fd_sc_hd__and2_1 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__nand3_1 (!A) | (!B) | (!C)
.model d_lut_sky130_fd_sc_hd__nand3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11111110")
* sky130_fd_sc_hd__and3b_1 (!A_N&B&C)
.model d_lut_sky130_fd_sc_hd__and3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000010")
* sky130_fd_sc_hd__and4_1 (A&B&C&D)
.model d_lut_sky130_fd_sc_hd__and4_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000001")
* sky130_fd_sc_hd__a21o_1 (A1&A2) | (B1)
.model d_lut_sky130_fd_sc_hd__a21o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00011111")
* sky130_fd_sc_hd__clkbuf_1 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__dlymetal6s2s_1 (A)
.model d_lut_sky130_fd_sc_hd__dlymetal6s2s_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__conb_1 1
* sky130_fd_sc_hd__a211o_1 (A1&A2) | (B1) | (C1)
.model d_lut_sky130_fd_sc_hd__a211o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001111111111111")
* sky130_fd_sc_hd__buf_1 (A)
.model d_lut_sky130_fd_sc_hd__buf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__nor2_2 (!A&!B)
.model d_lut_sky130_fd_sc_hd__nor2_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1000")
* sky130_fd_sc_hd__dfrtp_4 IQ
* sky130_fd_sc_hd__and4_2 (A&B&C&D)
.model d_lut_sky130_fd_sc_hd__and4_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000001")
* sky130_fd_sc_hd__diode_2 (no function)
.end

magic
tech sky130A
timestamp 1712352531
<< pwell >>
rect -856 -379 856 379
<< mvnmos >>
rect -742 -250 -682 250
rect -653 -250 -593 250
rect -564 -250 -504 250
rect -475 -250 -415 250
rect -386 -250 -326 250
rect -297 -250 -237 250
rect -208 -250 -148 250
rect -119 -250 -59 250
rect -30 -250 30 250
rect 59 -250 119 250
rect 148 -250 208 250
rect 237 -250 297 250
rect 326 -250 386 250
rect 415 -250 475 250
rect 504 -250 564 250
rect 593 -250 653 250
rect 682 -250 742 250
<< mvndiff >>
rect -771 244 -742 250
rect -771 -244 -765 244
rect -748 -244 -742 244
rect -771 -250 -742 -244
rect -682 244 -653 250
rect -682 -244 -676 244
rect -659 -244 -653 244
rect -682 -250 -653 -244
rect -593 244 -564 250
rect -593 -244 -587 244
rect -570 -244 -564 244
rect -593 -250 -564 -244
rect -504 244 -475 250
rect -504 -244 -498 244
rect -481 -244 -475 244
rect -504 -250 -475 -244
rect -415 244 -386 250
rect -415 -244 -409 244
rect -392 -244 -386 244
rect -415 -250 -386 -244
rect -326 244 -297 250
rect -326 -244 -320 244
rect -303 -244 -297 244
rect -326 -250 -297 -244
rect -237 244 -208 250
rect -237 -244 -231 244
rect -214 -244 -208 244
rect -237 -250 -208 -244
rect -148 244 -119 250
rect -148 -244 -142 244
rect -125 -244 -119 244
rect -148 -250 -119 -244
rect -59 244 -30 250
rect -59 -244 -53 244
rect -36 -244 -30 244
rect -59 -250 -30 -244
rect 30 244 59 250
rect 30 -244 36 244
rect 53 -244 59 244
rect 30 -250 59 -244
rect 119 244 148 250
rect 119 -244 125 244
rect 142 -244 148 244
rect 119 -250 148 -244
rect 208 244 237 250
rect 208 -244 214 244
rect 231 -244 237 244
rect 208 -250 237 -244
rect 297 244 326 250
rect 297 -244 303 244
rect 320 -244 326 244
rect 297 -250 326 -244
rect 386 244 415 250
rect 386 -244 392 244
rect 409 -244 415 244
rect 386 -250 415 -244
rect 475 244 504 250
rect 475 -244 481 244
rect 498 -244 504 244
rect 475 -250 504 -244
rect 564 244 593 250
rect 564 -244 570 244
rect 587 -244 593 244
rect 564 -250 593 -244
rect 653 244 682 250
rect 653 -244 659 244
rect 676 -244 682 244
rect 653 -250 682 -244
rect 742 244 771 250
rect 742 -244 748 244
rect 765 -244 771 244
rect 742 -250 771 -244
<< mvndiffc >>
rect -765 -244 -748 244
rect -676 -244 -659 244
rect -587 -244 -570 244
rect -498 -244 -481 244
rect -409 -244 -392 244
rect -320 -244 -303 244
rect -231 -244 -214 244
rect -142 -244 -125 244
rect -53 -244 -36 244
rect 36 -244 53 244
rect 125 -244 142 244
rect 214 -244 231 244
rect 303 -244 320 244
rect 392 -244 409 244
rect 481 -244 498 244
rect 570 -244 587 244
rect 659 -244 676 244
rect 748 -244 765 244
<< mvpsubdiff >>
rect -838 355 838 361
rect -838 338 -784 355
rect 784 338 838 355
rect -838 332 838 338
rect -838 307 -809 332
rect -838 -307 -832 307
rect -815 -307 -809 307
rect 809 307 838 332
rect -838 -332 -809 -307
rect 809 -307 815 307
rect 832 -307 838 307
rect 809 -332 838 -307
rect -838 -338 838 -332
rect -838 -355 -784 -338
rect 784 -355 838 -338
rect -838 -361 838 -355
<< mvpsubdiffcont >>
rect -784 338 784 355
rect -832 -307 -815 307
rect 815 -307 832 307
rect -784 -355 784 -338
<< poly >>
rect -742 286 -682 294
rect -742 269 -734 286
rect -690 269 -682 286
rect -742 250 -682 269
rect -653 286 -593 294
rect -653 269 -645 286
rect -601 269 -593 286
rect -653 250 -593 269
rect -564 286 -504 294
rect -564 269 -556 286
rect -512 269 -504 286
rect -564 250 -504 269
rect -475 286 -415 294
rect -475 269 -467 286
rect -423 269 -415 286
rect -475 250 -415 269
rect -386 286 -326 294
rect -386 269 -378 286
rect -334 269 -326 286
rect -386 250 -326 269
rect -297 286 -237 294
rect -297 269 -289 286
rect -245 269 -237 286
rect -297 250 -237 269
rect -208 286 -148 294
rect -208 269 -200 286
rect -156 269 -148 286
rect -208 250 -148 269
rect -119 286 -59 294
rect -119 269 -111 286
rect -67 269 -59 286
rect -119 250 -59 269
rect -30 286 30 294
rect -30 269 -22 286
rect 22 269 30 286
rect -30 250 30 269
rect 59 286 119 294
rect 59 269 67 286
rect 111 269 119 286
rect 59 250 119 269
rect 148 286 208 294
rect 148 269 156 286
rect 200 269 208 286
rect 148 250 208 269
rect 237 286 297 294
rect 237 269 245 286
rect 289 269 297 286
rect 237 250 297 269
rect 326 286 386 294
rect 326 269 334 286
rect 378 269 386 286
rect 326 250 386 269
rect 415 286 475 294
rect 415 269 423 286
rect 467 269 475 286
rect 415 250 475 269
rect 504 286 564 294
rect 504 269 512 286
rect 556 269 564 286
rect 504 250 564 269
rect 593 286 653 294
rect 593 269 601 286
rect 645 269 653 286
rect 593 250 653 269
rect 682 286 742 294
rect 682 269 690 286
rect 734 269 742 286
rect 682 250 742 269
rect -742 -269 -682 -250
rect -742 -286 -734 -269
rect -690 -286 -682 -269
rect -742 -294 -682 -286
rect -653 -269 -593 -250
rect -653 -286 -645 -269
rect -601 -286 -593 -269
rect -653 -294 -593 -286
rect -564 -269 -504 -250
rect -564 -286 -556 -269
rect -512 -286 -504 -269
rect -564 -294 -504 -286
rect -475 -269 -415 -250
rect -475 -286 -467 -269
rect -423 -286 -415 -269
rect -475 -294 -415 -286
rect -386 -269 -326 -250
rect -386 -286 -378 -269
rect -334 -286 -326 -269
rect -386 -294 -326 -286
rect -297 -269 -237 -250
rect -297 -286 -289 -269
rect -245 -286 -237 -269
rect -297 -294 -237 -286
rect -208 -269 -148 -250
rect -208 -286 -200 -269
rect -156 -286 -148 -269
rect -208 -294 -148 -286
rect -119 -269 -59 -250
rect -119 -286 -111 -269
rect -67 -286 -59 -269
rect -119 -294 -59 -286
rect -30 -269 30 -250
rect -30 -286 -22 -269
rect 22 -286 30 -269
rect -30 -294 30 -286
rect 59 -269 119 -250
rect 59 -286 67 -269
rect 111 -286 119 -269
rect 59 -294 119 -286
rect 148 -269 208 -250
rect 148 -286 156 -269
rect 200 -286 208 -269
rect 148 -294 208 -286
rect 237 -269 297 -250
rect 237 -286 245 -269
rect 289 -286 297 -269
rect 237 -294 297 -286
rect 326 -269 386 -250
rect 326 -286 334 -269
rect 378 -286 386 -269
rect 326 -294 386 -286
rect 415 -269 475 -250
rect 415 -286 423 -269
rect 467 -286 475 -269
rect 415 -294 475 -286
rect 504 -269 564 -250
rect 504 -286 512 -269
rect 556 -286 564 -269
rect 504 -294 564 -286
rect 593 -269 653 -250
rect 593 -286 601 -269
rect 645 -286 653 -269
rect 593 -294 653 -286
rect 682 -269 742 -250
rect 682 -286 690 -269
rect 734 -286 742 -269
rect 682 -294 742 -286
<< polycont >>
rect -734 269 -690 286
rect -645 269 -601 286
rect -556 269 -512 286
rect -467 269 -423 286
rect -378 269 -334 286
rect -289 269 -245 286
rect -200 269 -156 286
rect -111 269 -67 286
rect -22 269 22 286
rect 67 269 111 286
rect 156 269 200 286
rect 245 269 289 286
rect 334 269 378 286
rect 423 269 467 286
rect 512 269 556 286
rect 601 269 645 286
rect 690 269 734 286
rect -734 -286 -690 -269
rect -645 -286 -601 -269
rect -556 -286 -512 -269
rect -467 -286 -423 -269
rect -378 -286 -334 -269
rect -289 -286 -245 -269
rect -200 -286 -156 -269
rect -111 -286 -67 -269
rect -22 -286 22 -269
rect 67 -286 111 -269
rect 156 -286 200 -269
rect 245 -286 289 -269
rect 334 -286 378 -269
rect 423 -286 467 -269
rect 512 -286 556 -269
rect 601 -286 645 -269
rect 690 -286 734 -269
<< locali >>
rect -832 338 -784 355
rect 784 338 832 355
rect -832 307 -815 338
rect 815 307 832 338
rect -742 269 -734 286
rect -690 269 -682 286
rect -653 269 -645 286
rect -601 269 -593 286
rect -564 269 -556 286
rect -512 269 -504 286
rect -475 269 -467 286
rect -423 269 -415 286
rect -386 269 -378 286
rect -334 269 -326 286
rect -297 269 -289 286
rect -245 269 -237 286
rect -208 269 -200 286
rect -156 269 -148 286
rect -119 269 -111 286
rect -67 269 -59 286
rect -30 269 -22 286
rect 22 269 30 286
rect 59 269 67 286
rect 111 269 119 286
rect 148 269 156 286
rect 200 269 208 286
rect 237 269 245 286
rect 289 269 297 286
rect 326 269 334 286
rect 378 269 386 286
rect 415 269 423 286
rect 467 269 475 286
rect 504 269 512 286
rect 556 269 564 286
rect 593 269 601 286
rect 645 269 653 286
rect 682 269 690 286
rect 734 269 742 286
rect -765 244 -748 252
rect -765 -252 -748 -244
rect -676 244 -659 252
rect -676 -252 -659 -244
rect -587 244 -570 252
rect -587 -252 -570 -244
rect -498 244 -481 252
rect -498 -252 -481 -244
rect -409 244 -392 252
rect -409 -252 -392 -244
rect -320 244 -303 252
rect -320 -252 -303 -244
rect -231 244 -214 252
rect -231 -252 -214 -244
rect -142 244 -125 252
rect -142 -252 -125 -244
rect -53 244 -36 252
rect -53 -252 -36 -244
rect 36 244 53 252
rect 36 -252 53 -244
rect 125 244 142 252
rect 125 -252 142 -244
rect 214 244 231 252
rect 214 -252 231 -244
rect 303 244 320 252
rect 303 -252 320 -244
rect 392 244 409 252
rect 392 -252 409 -244
rect 481 244 498 252
rect 481 -252 498 -244
rect 570 244 587 252
rect 570 -252 587 -244
rect 659 244 676 252
rect 659 -252 676 -244
rect 748 244 765 252
rect 748 -252 765 -244
rect -742 -286 -734 -269
rect -690 -286 -682 -269
rect -653 -286 -645 -269
rect -601 -286 -593 -269
rect -564 -286 -556 -269
rect -512 -286 -504 -269
rect -475 -286 -467 -269
rect -423 -286 -415 -269
rect -386 -286 -378 -269
rect -334 -286 -326 -269
rect -297 -286 -289 -269
rect -245 -286 -237 -269
rect -208 -286 -200 -269
rect -156 -286 -148 -269
rect -119 -286 -111 -269
rect -67 -286 -59 -269
rect -30 -286 -22 -269
rect 22 -286 30 -269
rect 59 -286 67 -269
rect 111 -286 119 -269
rect 148 -286 156 -269
rect 200 -286 208 -269
rect 237 -286 245 -269
rect 289 -286 297 -269
rect 326 -286 334 -269
rect 378 -286 386 -269
rect 415 -286 423 -269
rect 467 -286 475 -269
rect 504 -286 512 -269
rect 556 -286 564 -269
rect 593 -286 601 -269
rect 645 -286 653 -269
rect 682 -286 690 -269
rect 734 -286 742 -269
rect -832 -338 -815 -307
rect 815 -338 832 -307
rect -832 -355 -784 -338
rect 784 -355 832 -338
<< viali >>
rect -734 269 -690 286
rect -645 269 -601 286
rect -556 269 -512 286
rect -467 269 -423 286
rect -378 269 -334 286
rect -289 269 -245 286
rect -200 269 -156 286
rect -111 269 -67 286
rect -22 269 22 286
rect 67 269 111 286
rect 156 269 200 286
rect 245 269 289 286
rect 334 269 378 286
rect 423 269 467 286
rect 512 269 556 286
rect 601 269 645 286
rect 690 269 734 286
rect -765 -244 -748 244
rect -676 -244 -659 244
rect -587 -244 -570 244
rect -498 -244 -481 244
rect -409 -244 -392 244
rect -320 -244 -303 244
rect -231 -244 -214 244
rect -142 -244 -125 244
rect -53 -244 -36 244
rect 36 -244 53 244
rect 125 -244 142 244
rect 214 -244 231 244
rect 303 -244 320 244
rect 392 -244 409 244
rect 481 -244 498 244
rect 570 -244 587 244
rect 659 -244 676 244
rect 748 -244 765 244
rect -734 -286 -690 -269
rect -645 -286 -601 -269
rect -556 -286 -512 -269
rect -467 -286 -423 -269
rect -378 -286 -334 -269
rect -289 -286 -245 -269
rect -200 -286 -156 -269
rect -111 -286 -67 -269
rect -22 -286 22 -269
rect 67 -286 111 -269
rect 156 -286 200 -269
rect 245 -286 289 -269
rect 334 -286 378 -269
rect 423 -286 467 -269
rect 512 -286 556 -269
rect 601 -286 645 -269
rect 690 -286 734 -269
<< metal1 >>
rect -740 286 -684 289
rect -740 269 -734 286
rect -690 269 -684 286
rect -740 266 -684 269
rect -651 286 -595 289
rect -651 269 -645 286
rect -601 269 -595 286
rect -651 266 -595 269
rect -562 286 -506 289
rect -562 269 -556 286
rect -512 269 -506 286
rect -562 266 -506 269
rect -473 286 -417 289
rect -473 269 -467 286
rect -423 269 -417 286
rect -473 266 -417 269
rect -384 286 -328 289
rect -384 269 -378 286
rect -334 269 -328 286
rect -384 266 -328 269
rect -295 286 -239 289
rect -295 269 -289 286
rect -245 269 -239 286
rect -295 266 -239 269
rect -206 286 -150 289
rect -206 269 -200 286
rect -156 269 -150 286
rect -206 266 -150 269
rect -117 286 -61 289
rect -117 269 -111 286
rect -67 269 -61 286
rect -117 266 -61 269
rect -28 286 28 289
rect -28 269 -22 286
rect 22 269 28 286
rect -28 266 28 269
rect 61 286 117 289
rect 61 269 67 286
rect 111 269 117 286
rect 61 266 117 269
rect 150 286 206 289
rect 150 269 156 286
rect 200 269 206 286
rect 150 266 206 269
rect 239 286 295 289
rect 239 269 245 286
rect 289 269 295 286
rect 239 266 295 269
rect 328 286 384 289
rect 328 269 334 286
rect 378 269 384 286
rect 328 266 384 269
rect 417 286 473 289
rect 417 269 423 286
rect 467 269 473 286
rect 417 266 473 269
rect 506 286 562 289
rect 506 269 512 286
rect 556 269 562 286
rect 506 266 562 269
rect 595 286 651 289
rect 595 269 601 286
rect 645 269 651 286
rect 595 266 651 269
rect 684 286 740 289
rect 684 269 690 286
rect 734 269 740 286
rect 684 266 740 269
rect -768 244 -745 250
rect -768 -244 -765 244
rect -748 -244 -745 244
rect -768 -250 -745 -244
rect -679 244 -656 250
rect -679 -244 -676 244
rect -659 -244 -656 244
rect -679 -250 -656 -244
rect -590 244 -567 250
rect -590 -244 -587 244
rect -570 -244 -567 244
rect -590 -250 -567 -244
rect -501 244 -478 250
rect -501 -244 -498 244
rect -481 -244 -478 244
rect -501 -250 -478 -244
rect -412 244 -389 250
rect -412 -244 -409 244
rect -392 -244 -389 244
rect -412 -250 -389 -244
rect -323 244 -300 250
rect -323 -244 -320 244
rect -303 -244 -300 244
rect -323 -250 -300 -244
rect -234 244 -211 250
rect -234 -244 -231 244
rect -214 -244 -211 244
rect -234 -250 -211 -244
rect -145 244 -122 250
rect -145 -244 -142 244
rect -125 -244 -122 244
rect -145 -250 -122 -244
rect -56 244 -33 250
rect -56 -244 -53 244
rect -36 -244 -33 244
rect -56 -250 -33 -244
rect 33 244 56 250
rect 33 -244 36 244
rect 53 -244 56 244
rect 33 -250 56 -244
rect 122 244 145 250
rect 122 -244 125 244
rect 142 -244 145 244
rect 122 -250 145 -244
rect 211 244 234 250
rect 211 -244 214 244
rect 231 -244 234 244
rect 211 -250 234 -244
rect 300 244 323 250
rect 300 -244 303 244
rect 320 -244 323 244
rect 300 -250 323 -244
rect 389 244 412 250
rect 389 -244 392 244
rect 409 -244 412 244
rect 389 -250 412 -244
rect 478 244 501 250
rect 478 -244 481 244
rect 498 -244 501 244
rect 478 -250 501 -244
rect 567 244 590 250
rect 567 -244 570 244
rect 587 -244 590 244
rect 567 -250 590 -244
rect 656 244 679 250
rect 656 -244 659 244
rect 676 -244 679 244
rect 656 -250 679 -244
rect 745 244 768 250
rect 745 -244 748 244
rect 765 -244 768 244
rect 745 -250 768 -244
rect -740 -269 -684 -266
rect -740 -286 -734 -269
rect -690 -286 -684 -269
rect -740 -289 -684 -286
rect -651 -269 -595 -266
rect -651 -286 -645 -269
rect -601 -286 -595 -269
rect -651 -289 -595 -286
rect -562 -269 -506 -266
rect -562 -286 -556 -269
rect -512 -286 -506 -269
rect -562 -289 -506 -286
rect -473 -269 -417 -266
rect -473 -286 -467 -269
rect -423 -286 -417 -269
rect -473 -289 -417 -286
rect -384 -269 -328 -266
rect -384 -286 -378 -269
rect -334 -286 -328 -269
rect -384 -289 -328 -286
rect -295 -269 -239 -266
rect -295 -286 -289 -269
rect -245 -286 -239 -269
rect -295 -289 -239 -286
rect -206 -269 -150 -266
rect -206 -286 -200 -269
rect -156 -286 -150 -269
rect -206 -289 -150 -286
rect -117 -269 -61 -266
rect -117 -286 -111 -269
rect -67 -286 -61 -269
rect -117 -289 -61 -286
rect -28 -269 28 -266
rect -28 -286 -22 -269
rect 22 -286 28 -269
rect -28 -289 28 -286
rect 61 -269 117 -266
rect 61 -286 67 -269
rect 111 -286 117 -269
rect 61 -289 117 -286
rect 150 -269 206 -266
rect 150 -286 156 -269
rect 200 -286 206 -269
rect 150 -289 206 -286
rect 239 -269 295 -266
rect 239 -286 245 -269
rect 289 -286 295 -269
rect 239 -289 295 -286
rect 328 -269 384 -266
rect 328 -286 334 -269
rect 378 -286 384 -269
rect 328 -289 384 -286
rect 417 -269 473 -266
rect 417 -286 423 -269
rect 467 -286 473 -269
rect 417 -289 473 -286
rect 506 -269 562 -266
rect 506 -286 512 -269
rect 556 -286 562 -269
rect 506 -289 562 -286
rect 595 -269 651 -266
rect 595 -286 601 -269
rect 645 -286 651 -269
rect 595 -289 651 -286
rect 684 -269 740 -266
rect 684 -286 690 -269
rect 734 -286 740 -269
rect 684 -289 740 -286
<< properties >>
string FIXED_BBOX -823 -346 823 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 17 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712930986
<< pwell >>
rect -5173 -505 5173 505
<< mvnmos >>
rect -4945 47 -3345 247
rect -3287 47 -1687 247
rect -1629 47 -29 247
rect 29 47 1629 247
rect 1687 47 3287 247
rect 3345 47 4945 247
rect -4945 -309 -3345 -109
rect -3287 -309 -1687 -109
rect -1629 -309 -29 -109
rect 29 -309 1629 -109
rect 1687 -309 3287 -109
rect 3345 -309 4945 -109
<< mvndiff >>
rect -5003 235 -4945 247
rect -5003 59 -4991 235
rect -4957 59 -4945 235
rect -5003 47 -4945 59
rect -3345 235 -3287 247
rect -3345 59 -3333 235
rect -3299 59 -3287 235
rect -3345 47 -3287 59
rect -1687 235 -1629 247
rect -1687 59 -1675 235
rect -1641 59 -1629 235
rect -1687 47 -1629 59
rect -29 235 29 247
rect -29 59 -17 235
rect 17 59 29 235
rect -29 47 29 59
rect 1629 235 1687 247
rect 1629 59 1641 235
rect 1675 59 1687 235
rect 1629 47 1687 59
rect 3287 235 3345 247
rect 3287 59 3299 235
rect 3333 59 3345 235
rect 3287 47 3345 59
rect 4945 235 5003 247
rect 4945 59 4957 235
rect 4991 59 5003 235
rect 4945 47 5003 59
rect -5003 -121 -4945 -109
rect -5003 -297 -4991 -121
rect -4957 -297 -4945 -121
rect -5003 -309 -4945 -297
rect -3345 -121 -3287 -109
rect -3345 -297 -3333 -121
rect -3299 -297 -3287 -121
rect -3345 -309 -3287 -297
rect -1687 -121 -1629 -109
rect -1687 -297 -1675 -121
rect -1641 -297 -1629 -121
rect -1687 -309 -1629 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 1629 -121 1687 -109
rect 1629 -297 1641 -121
rect 1675 -297 1687 -121
rect 1629 -309 1687 -297
rect 3287 -121 3345 -109
rect 3287 -297 3299 -121
rect 3333 -297 3345 -121
rect 3287 -309 3345 -297
rect 4945 -121 5003 -109
rect 4945 -297 4957 -121
rect 4991 -297 5003 -121
rect 4945 -309 5003 -297
<< mvndiffc >>
rect -4991 59 -4957 235
rect -3333 59 -3299 235
rect -1675 59 -1641 235
rect -17 59 17 235
rect 1641 59 1675 235
rect 3299 59 3333 235
rect 4957 59 4991 235
rect -4991 -297 -4957 -121
rect -3333 -297 -3299 -121
rect -1675 -297 -1641 -121
rect -17 -297 17 -121
rect 1641 -297 1675 -121
rect 3299 -297 3333 -121
rect 4957 -297 4991 -121
<< mvpsubdiff >>
rect -5137 457 5137 469
rect -5137 423 -5029 457
rect 5029 423 5137 457
rect -5137 411 5137 423
rect -5137 361 -5079 411
rect -5137 -361 -5125 361
rect -5091 -361 -5079 361
rect 5079 361 5137 411
rect -5137 -411 -5079 -361
rect 5079 -361 5091 361
rect 5125 -361 5137 361
rect 5079 -411 5137 -361
rect -5137 -423 5137 -411
rect -5137 -457 -5029 -423
rect 5029 -457 5137 -423
rect -5137 -469 5137 -457
<< mvpsubdiffcont >>
rect -5029 423 5029 457
rect -5125 -361 -5091 361
rect 5091 -361 5125 361
rect -5029 -457 5029 -423
<< poly >>
rect -4945 319 -3345 335
rect -4945 285 -4929 319
rect -3361 285 -3345 319
rect -4945 247 -3345 285
rect -3287 319 -1687 335
rect -3287 285 -3271 319
rect -1703 285 -1687 319
rect -3287 247 -1687 285
rect -1629 319 -29 335
rect -1629 285 -1613 319
rect -45 285 -29 319
rect -1629 247 -29 285
rect 29 319 1629 335
rect 29 285 45 319
rect 1613 285 1629 319
rect 29 247 1629 285
rect 1687 319 3287 335
rect 1687 285 1703 319
rect 3271 285 3287 319
rect 1687 247 3287 285
rect 3345 319 4945 335
rect 3345 285 3361 319
rect 4929 285 4945 319
rect 3345 247 4945 285
rect -4945 21 -3345 47
rect -3287 21 -1687 47
rect -1629 21 -29 47
rect 29 21 1629 47
rect 1687 21 3287 47
rect 3345 21 4945 47
rect -4945 -37 -3345 -21
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -4945 -109 -3345 -71
rect -3287 -37 -1687 -21
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -3287 -109 -1687 -71
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -109 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -109 1629 -71
rect 1687 -37 3287 -21
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 1687 -109 3287 -71
rect 3345 -37 4945 -21
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 3345 -109 4945 -71
rect -4945 -335 -3345 -309
rect -3287 -335 -1687 -309
rect -1629 -335 -29 -309
rect 29 -335 1629 -309
rect 1687 -335 3287 -309
rect 3345 -335 4945 -309
<< polycont >>
rect -4929 285 -3361 319
rect -3271 285 -1703 319
rect -1613 285 -45 319
rect 45 285 1613 319
rect 1703 285 3271 319
rect 3361 285 4929 319
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
<< locali >>
rect -5125 423 -5029 457
rect 5029 423 5125 457
rect -5125 361 -5091 423
rect 5091 361 5125 423
rect -4945 285 -4929 319
rect -3361 285 -3345 319
rect -3287 285 -3271 319
rect -1703 285 -1687 319
rect -1629 285 -1613 319
rect -45 285 -29 319
rect 29 285 45 319
rect 1613 285 1629 319
rect 1687 285 1703 319
rect 3271 285 3287 319
rect 3345 285 3361 319
rect 4929 285 4945 319
rect -4991 235 -4957 251
rect -4991 43 -4957 59
rect -3333 235 -3299 251
rect -3333 43 -3299 59
rect -1675 235 -1641 251
rect -1675 43 -1641 59
rect -17 235 17 251
rect -17 43 17 59
rect 1641 235 1675 251
rect 1641 43 1675 59
rect 3299 235 3333 251
rect 3299 43 3333 59
rect 4957 235 4991 251
rect 4957 43 4991 59
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect -4991 -121 -4957 -105
rect -4991 -313 -4957 -297
rect -3333 -121 -3299 -105
rect -3333 -313 -3299 -297
rect -1675 -121 -1641 -105
rect -1675 -313 -1641 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 1641 -121 1675 -105
rect 1641 -313 1675 -297
rect 3299 -121 3333 -105
rect 3299 -313 3333 -297
rect 4957 -121 4991 -105
rect 4957 -313 4991 -297
rect -5125 -423 -5091 -361
rect 5091 -423 5125 -361
rect -5125 -457 -5029 -423
rect 5029 -457 5125 -423
<< viali >>
rect -4929 285 -3361 319
rect -3271 285 -1703 319
rect -1613 285 -45 319
rect 45 285 1613 319
rect 1703 285 3271 319
rect 3361 285 4929 319
rect -4991 59 -4957 235
rect -3333 59 -3299 235
rect -1675 59 -1641 235
rect -17 59 17 235
rect 1641 59 1675 235
rect 3299 59 3333 235
rect 4957 59 4991 235
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect -4991 -297 -4957 -121
rect -3333 -297 -3299 -121
rect -1675 -297 -1641 -121
rect -17 -297 17 -121
rect 1641 -297 1675 -121
rect 3299 -297 3333 -121
rect 4957 -297 4991 -121
<< metal1 >>
rect -4941 319 -3349 325
rect -4941 285 -4929 319
rect -3361 285 -3349 319
rect -4941 279 -3349 285
rect -3283 319 -1691 325
rect -3283 285 -3271 319
rect -1703 285 -1691 319
rect -3283 279 -1691 285
rect -1625 319 -33 325
rect -1625 285 -1613 319
rect -45 285 -33 319
rect -1625 279 -33 285
rect 33 319 1625 325
rect 33 285 45 319
rect 1613 285 1625 319
rect 33 279 1625 285
rect 1691 319 3283 325
rect 1691 285 1703 319
rect 3271 285 3283 319
rect 1691 279 3283 285
rect 3349 319 4941 325
rect 3349 285 3361 319
rect 4929 285 4941 319
rect 3349 279 4941 285
rect -4997 235 -4951 247
rect -4997 59 -4991 235
rect -4957 59 -4951 235
rect -4997 47 -4951 59
rect -3339 235 -3293 247
rect -3339 59 -3333 235
rect -3299 59 -3293 235
rect -3339 47 -3293 59
rect -1681 235 -1635 247
rect -1681 59 -1675 235
rect -1641 59 -1635 235
rect -1681 47 -1635 59
rect -23 235 23 247
rect -23 59 -17 235
rect 17 59 23 235
rect -23 47 23 59
rect 1635 235 1681 247
rect 1635 59 1641 235
rect 1675 59 1681 235
rect 1635 47 1681 59
rect 3293 235 3339 247
rect 3293 59 3299 235
rect 3333 59 3339 235
rect 3293 47 3339 59
rect 4951 235 4997 247
rect 4951 59 4957 235
rect 4991 59 4997 235
rect 4951 47 4997 59
rect -4941 -37 -3349 -31
rect -4941 -71 -4929 -37
rect -3361 -71 -3349 -37
rect -4941 -77 -3349 -71
rect -3283 -37 -1691 -31
rect -3283 -71 -3271 -37
rect -1703 -71 -1691 -37
rect -3283 -77 -1691 -71
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect 1691 -37 3283 -31
rect 1691 -71 1703 -37
rect 3271 -71 3283 -37
rect 1691 -77 3283 -71
rect 3349 -37 4941 -31
rect 3349 -71 3361 -37
rect 4929 -71 4941 -37
rect 3349 -77 4941 -71
rect -4997 -121 -4951 -109
rect -4997 -297 -4991 -121
rect -4957 -297 -4951 -121
rect -4997 -309 -4951 -297
rect -3339 -121 -3293 -109
rect -3339 -297 -3333 -121
rect -3299 -297 -3293 -121
rect -3339 -309 -3293 -297
rect -1681 -121 -1635 -109
rect -1681 -297 -1675 -121
rect -1641 -297 -1635 -121
rect -1681 -309 -1635 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 1635 -121 1681 -109
rect 1635 -297 1641 -121
rect 1675 -297 1681 -121
rect 1635 -309 1681 -297
rect 3293 -121 3339 -109
rect 3293 -297 3299 -121
rect 3333 -297 3339 -121
rect 3293 -309 3339 -297
rect 4951 -121 4997 -109
rect 4951 -297 4957 -121
rect 4991 -297 4997 -121
rect 4951 -309 4997 -297
<< properties >>
string FIXED_BBOX -5108 -440 5108 440
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 8 m 2 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

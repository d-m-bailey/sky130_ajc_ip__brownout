* NGSPICE file created from sky130_ef_sc_hd__fill_8.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__fill_8 abstract view
.subckt sky130_ef_sc_hd__fill_8 VPWR VGND VPB VNB
.ends


* NGSPICE file created from brownout_dig.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt brownout_dig VGND VPWR brout_filt ena force_rc_osc force_short_oneshot osc_ck
+ osc_ck_256 osc_ena otrip[0] otrip[1] otrip[2] otrip_decoded[0] otrip_decoded[1]
+ otrip_decoded[2] otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6]
+ otrip_decoded[7] out_unbuf timed_out vtrip[0] vtrip[1] vtrip[2] vtrip_decoded[0]
+ vtrip_decoded[1] vtrip_decoded[2] vtrip_decoded[3] vtrip_decoded[4] vtrip_decoded[5]
+ vtrip_decoded[6] vtrip_decoded[7]
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_131_ cnt\[10\] net31 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_114_ _033_ _038_ net32 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput20 net20 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ cnt\[9\] cnt\[8\] _067_ net4 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_3__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_113_ _063_ _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR out_unbuf sky130_fd_sc_hd__buf_2
XFILLER_0_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_189_ clknet_2_2__leaf_osc_ck _005_ net37 VGND VGND VPWR VPWR cnt_ck_256\[5\] sky130_fd_sc_hd__dfrtp_1
X_112_ cnt\[1\] cnt\[0\] cnt\[2\] cnt\[3\] VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold10 cnt_ck_256\[1\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput22 net22 VGND VGND VPWR VPWR timed_out sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR osc_ck_256 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_188_ clknet_2_2__leaf_osc_ck _004_ net37 VGND VGND VPWR VPWR cnt_ck_256\[4\] sky130_fd_sc_hd__dfrtp_1
X_111_ _033_ _036_ net43 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold11 _001_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR vtrip_decoded[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_187_ clknet_2_2__leaf_osc_ck _003_ net37 VGND VGND VPWR VPWR cnt_ck_256\[3\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_8_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ cnt\[2\] _062_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__xor2_1
Xhold12 cnt_ck_256\[0\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput24 net24 VGND VGND VPWR VPWR vtrip_decoded[1] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_186_ clknet_2_3__leaf_osc_ck _002_ net37 VGND VGND VPWR VPWR cnt_ck_256\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ clknet_2_3__leaf_osc_ck _008_ net34 VGND VGND VPWR VPWR cnt\[1\] sky130_fd_sc_hd__dfstp_1
Xhold13 cnt_ck_256\[5\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_11_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput25 net25 VGND VGND VPWR VPWR vtrip_decoded[2] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_3_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ clknet_2_3__leaf_osc_ck net47 net37 VGND VGND VPWR VPWR cnt_ck_256\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_168_ clknet_2_3__leaf_osc_ck _007_ net34 VGND VGND VPWR VPWR cnt\[0\] sky130_fd_sc_hd__dfstp_1
X_099_ cnt_ck_256\[5\] cnt_ck_256\[4\] _027_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and3_1
Xhold14 _030_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR vtrip_decoded[3] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_184_ clknet_2_3__leaf_osc_ck _000_ net37 VGND VGND VPWR VPWR cnt_ck_256\[0\] sky130_fd_sc_hd__dfrtp_1
X_098_ net51 _027_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__xor2_1
X_167_ net7 net6 net5 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__nor3b_1
XFILLER_0_11_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 cnt_ck_256\[4\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR vtrip_decoded[4] sky130_fd_sc_hd__buf_2
XFILLER_0_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ clknet_2_0__leaf_osc_ck _022_ net33 VGND VGND VPWR VPWR cnt\[15\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_9_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_097_ _027_ _028_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nor2_1
X_166_ net7 net5 net6 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_19_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 cnt_ck_256\[2\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
X_149_ net45 _031_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VPWR VPWR vtrip_decoded[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ clknet_2_0__leaf_osc_ck _021_ net33 VGND VGND VPWR VPWR cnt\[14\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_0_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_165_ _073_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__inv_2
X_096_ net53 _025_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold17 cnt_ck_256\[3\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
X_148_ _061_ _059_ _060_ _024_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_079_ net7 net5 net6 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and3_1
Xoutput29 net29 VGND VGND VPWR VPWR vtrip_decoded[6] sky130_fd_sc_hd__buf_2
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_2__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_2__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout31 _048_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_181_ clknet_2_1__leaf_osc_ck _020_ net33 VGND VGND VPWR VPWR cnt\[13\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ _061_ net22 VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__nand2_1
X_095_ cnt_ck_256\[3\] _025_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_147_ cnt\[15\] _071_ net31 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_078_ net5 net6 net7 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and3b_1
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ clknet_2_3__leaf_osc_ck _019_ net33 VGND VGND VPWR VPWR cnt\[12\] sky130_fd_sc_hd__dfstp_1
Xfanout32 brout_filt_retimed VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_163_ cnt\[9\] cnt\[8\] _067_ _072_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__and4_1
X_094_ _025_ _026_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ net6 net5 net7 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and3b_1
X_146_ _071_ net31 cnt\[15\] VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_129_ _033_ _047_ net32 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout33 net42 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
X_162_ cnt\[14\] cnt\[15\] _070_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__and3_1
X_093_ cnt_ck_256\[0\] net46 net52 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_7_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 brout_filt VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_145_ _061_ _057_ _058_ _024_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ net5 net6 net7 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__nor3b_1
XFILLER_0_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_128_ _068_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout34 net42 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
X_161_ cnt\[14\] _070_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ cnt_ck_256\[0\] cnt_ck_256\[1\] cnt_ck_256\[2\] VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and3_1
Xinput2 ena VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_075_ net7 net5 net6 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and3b_1
X_144_ _071_ net31 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197__36 VGND VGND VPWR VPWR net36 _197__36/LO sky130_fd_sc_hd__conb_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_127_ cnt\[8\] _067_ cnt\[9\] VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_10_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_160_ cnt\[11\] cnt\[10\] cnt\[13\] cnt\[12\] VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__and4_1
X_091_ cnt_ck_256\[0\] net46 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__xor2_1
Xinput3 force_rc_osc VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_143_ _070_ net31 cnt\[14\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__a21o_1
X_074_ net7 net5 net6 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
X_126_ _033_ _045_ net32 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ _033_ _035_ net43 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_090_ net2 _073_ brout_filt_ena_rsb net3 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__a211o_1
Xinput4 force_short_oneshot VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_142_ _055_ _056_ _024_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_125_ cnt\[8\] _067_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_108_ _062_ _034_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 otrip[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_141_ _070_ _048_ net32 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_124_ _033_ _044_ net32 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_14_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 otrip[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_2_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_140_ _069_ _048_ cnt\[13\] VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ cnt\[7\] _066_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__xnor2_1
X_106_ net44 _033_ net43 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 otrip[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_122_ _033_ _043_ net32 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 vtrip[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_2_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_105_ net4 net22 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 vtrip[0] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
X_198_ clknet_2_2__leaf_osc_ck net39 brout_filt_ena_rsb VGND VGND VPWR VPWR brout_filt_retime_rsb
+ sky130_fd_sc_hd__dfrtp_4
X_121_ _066_ _042_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_104_ _031_ _032_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 vtrip[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
X_197_ clknet_2_0__leaf_osc_ck net36 brout_filt_ena_rsb VGND VGND VPWR VPWR brout_filt_retime_rsb_stg1
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ cnt\[5\] cnt\[4\] _063_ cnt\[6\] VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_6_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ cnt_ck_256\[6\] _029_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 brout_filt_retime_rsb VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_14_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_196_ clknet_2_2__leaf_osc_ck net38 net37 VGND VGND VPWR VPWR brout_filt_retimed
+ sky130_fd_sc_hd__dfrtp_1
X_179_ clknet_2_2__leaf_osc_ck _018_ net33 VGND VGND VPWR VPWR cnt\[11\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
X_102_ cnt_ck_256\[6\] _029_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 brout_filt_retimed_stg1 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_195_ clknet_2_0__leaf_osc_ck net1 net37 VGND VGND VPWR VPWR brout_filt_retimed_stg1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_178_ clknet_2_2__leaf_osc_ck _017_ net33 VGND VGND VPWR VPWR cnt\[10\] sky130_fd_sc_hd__dfstp_1
X_101_ _029_ net50 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nor2_1
Xhold3 brout_filt_retime_rsb_stg1 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_194_ clknet_2_0__leaf_osc_ck net41 net2 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_177_ clknet_2_1__leaf_osc_ck _016_ net33 VGND VGND VPWR VPWR cnt\[9\] sky130_fd_sc_hd__dfstp_1
X_100_ cnt_ck_256\[4\] _027_ net49 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 cnt_rsb_stg1 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_193_ clknet_2_0__leaf_osc_ck net40 net2 VGND VGND VPWR VPWR cnt_rsb_stg2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_176_ clknet_2_1__leaf_osc_ck _015_ net33 VGND VGND VPWR VPWR cnt\[8\] sky130_fd_sc_hd__dfstp_1
X_159_ cnt\[11\] cnt\[10\] cnt\[12\] VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 cnt_rsb_stg2 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_192_ clknet_2_0__leaf_osc_ck net35 net2 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_175_ clknet_2_1__leaf_osc_ck _014_ net33 VGND VGND VPWR VPWR cnt\[7\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_1_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_158_ cnt\[9\] cnt\[8\] _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__and3_1
X_089_ net1 net2 VGND VGND VPWR VPWR brout_filt_ena_rsb sky130_fd_sc_hd__and2_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 cnt_rsb VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_191_ clknet_2_2__leaf_osc_ck _023_ net37 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
X_174_ clknet_2_1__leaf_osc_ck _013_ net33 VGND VGND VPWR VPWR cnt\[6\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_157_ cnt\[4\] cnt\[7\] _063_ _065_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__and4_1
X_088_ _061_ cnt\[15\] _068_ _071_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__and4_2
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 brout_filt_retimed VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ clknet_2_2__leaf_osc_ck _006_ net37 VGND VGND VPWR VPWR cnt_ck_256\[6\] sky130_fd_sc_hd__dfrtp_1
X_173_ clknet_2_1__leaf_osc_ck _012_ net34 VGND VGND VPWR VPWR cnt\[5\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_156_ cnt\[4\] _063_ _065_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__and3_1
X_087_ net10 net9 net8 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_17_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 cnt\[0\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_139_ _053_ _054_ _024_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ clknet_2_1__leaf_osc_ck _011_ net34 VGND VGND VPWR VPWR cnt\[4\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_5_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_086_ net8 net9 net10 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__and3b_1
X_155_ cnt\[5\] cnt\[6\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 net11 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
X_138_ _069_ net31 net32 VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_171_ clknet_2_3__leaf_osc_ck _010_ net34 VGND VGND VPWR VPWR cnt\[3\] sky130_fd_sc_hd__dfstp_1
X_085_ net9 net8 net10 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__and3b_1
X_154_ cnt\[4\] _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_137_ cnt\[11\] cnt\[10\] net31 cnt\[12\] VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ clknet_2_3__leaf_osc_ck _009_ net34 VGND VGND VPWR VPWR cnt\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ net9 net8 net10 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_8_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ cnt\[1\] cnt\[0\] cnt\[3\] cnt\[2\] VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__and4_1
X_136_ _061_ _051_ _052_ _024_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_119_ _033_ _041_ net32 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_192__35 VGND VGND VPWR VPWR net35 _192__35/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ net10 net9 net8 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__and3b_1
X_152_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ cnt\[11\] cnt\[10\] net31 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nand3_1
X_118_ cnt\[5\] _064_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 otrip[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_082_ net10 net8 net9 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__nor3b_1
X_151_ net32 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_134_ cnt\[10\] net31 cnt\[11\] VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__a21o_1
X_117_ _033_ _040_ net32 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_12_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_081_ net10 net9 net8 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_0_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_150_ net48 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_133_ _061_ _049_ _050_ _024_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_116_ _064_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_080_ net10 net9 net8 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__nor3_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_132_ cnt\[10\] net31 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_115_ cnt\[4\] _063_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_5_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput30 net30 VGND VGND VPWR VPWR vtrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends


magic
tech sky130A
magscale 1 2
timestamp 1712422266
<< nwell >>
rect -1194 -284 1194 284
<< pmos >>
rect -998 -64 -898 136
rect -840 -64 -740 136
rect -682 -64 -582 136
rect -524 -64 -424 136
rect -366 -64 -266 136
rect -208 -64 -108 136
rect -50 -64 50 136
rect 108 -64 208 136
rect 266 -64 366 136
rect 424 -64 524 136
rect 582 -64 682 136
rect 740 -64 840 136
rect 898 -64 998 136
<< pdiff >>
rect -1056 124 -998 136
rect -1056 -52 -1044 124
rect -1010 -52 -998 124
rect -1056 -64 -998 -52
rect -898 124 -840 136
rect -898 -52 -886 124
rect -852 -52 -840 124
rect -898 -64 -840 -52
rect -740 124 -682 136
rect -740 -52 -728 124
rect -694 -52 -682 124
rect -740 -64 -682 -52
rect -582 124 -524 136
rect -582 -52 -570 124
rect -536 -52 -524 124
rect -582 -64 -524 -52
rect -424 124 -366 136
rect -424 -52 -412 124
rect -378 -52 -366 124
rect -424 -64 -366 -52
rect -266 124 -208 136
rect -266 -52 -254 124
rect -220 -52 -208 124
rect -266 -64 -208 -52
rect -108 124 -50 136
rect -108 -52 -96 124
rect -62 -52 -50 124
rect -108 -64 -50 -52
rect 50 124 108 136
rect 50 -52 62 124
rect 96 -52 108 124
rect 50 -64 108 -52
rect 208 124 266 136
rect 208 -52 220 124
rect 254 -52 266 124
rect 208 -64 266 -52
rect 366 124 424 136
rect 366 -52 378 124
rect 412 -52 424 124
rect 366 -64 424 -52
rect 524 124 582 136
rect 524 -52 536 124
rect 570 -52 582 124
rect 524 -64 582 -52
rect 682 124 740 136
rect 682 -52 694 124
rect 728 -52 740 124
rect 682 -64 740 -52
rect 840 124 898 136
rect 840 -52 852 124
rect 886 -52 898 124
rect 840 -64 898 -52
rect 998 124 1056 136
rect 998 -52 1010 124
rect 1044 -52 1056 124
rect 998 -64 1056 -52
<< pdiffc >>
rect -1044 -52 -1010 124
rect -886 -52 -852 124
rect -728 -52 -694 124
rect -570 -52 -536 124
rect -412 -52 -378 124
rect -254 -52 -220 124
rect -96 -52 -62 124
rect 62 -52 96 124
rect 220 -52 254 124
rect 378 -52 412 124
rect 536 -52 570 124
rect 694 -52 728 124
rect 852 -52 886 124
rect 1010 -52 1044 124
<< nsubdiff >>
rect -1158 214 -1062 248
rect 1062 214 1158 248
rect -1158 151 -1124 214
rect 1124 151 1158 214
rect -1158 -214 -1124 -151
rect 1124 -214 1158 -151
rect -1158 -248 -1062 -214
rect 1062 -248 1158 -214
<< nsubdiffcont >>
rect -1062 214 1062 248
rect -1158 -151 -1124 151
rect 1124 -151 1158 151
rect -1062 -248 1062 -214
<< poly >>
rect -998 136 -898 162
rect -840 136 -740 162
rect -682 136 -582 162
rect -524 136 -424 162
rect -366 136 -266 162
rect -208 136 -108 162
rect -50 136 50 162
rect 108 136 208 162
rect 266 136 366 162
rect 424 136 524 162
rect 582 136 682 162
rect 740 136 840 162
rect 898 136 998 162
rect -998 -111 -898 -64
rect -998 -145 -982 -111
rect -914 -145 -898 -111
rect -998 -161 -898 -145
rect -840 -111 -740 -64
rect -840 -145 -824 -111
rect -756 -145 -740 -111
rect -840 -161 -740 -145
rect -682 -111 -582 -64
rect -682 -145 -666 -111
rect -598 -145 -582 -111
rect -682 -161 -582 -145
rect -524 -111 -424 -64
rect -524 -145 -508 -111
rect -440 -145 -424 -111
rect -524 -161 -424 -145
rect -366 -111 -266 -64
rect -366 -145 -350 -111
rect -282 -145 -266 -111
rect -366 -161 -266 -145
rect -208 -111 -108 -64
rect -208 -145 -192 -111
rect -124 -145 -108 -111
rect -208 -161 -108 -145
rect -50 -111 50 -64
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect -50 -161 50 -145
rect 108 -111 208 -64
rect 108 -145 124 -111
rect 192 -145 208 -111
rect 108 -161 208 -145
rect 266 -111 366 -64
rect 266 -145 282 -111
rect 350 -145 366 -111
rect 266 -161 366 -145
rect 424 -111 524 -64
rect 424 -145 440 -111
rect 508 -145 524 -111
rect 424 -161 524 -145
rect 582 -111 682 -64
rect 582 -145 598 -111
rect 666 -145 682 -111
rect 582 -161 682 -145
rect 740 -111 840 -64
rect 740 -145 756 -111
rect 824 -145 840 -111
rect 740 -161 840 -145
rect 898 -111 998 -64
rect 898 -145 914 -111
rect 982 -145 998 -111
rect 898 -161 998 -145
<< polycont >>
rect -982 -145 -914 -111
rect -824 -145 -756 -111
rect -666 -145 -598 -111
rect -508 -145 -440 -111
rect -350 -145 -282 -111
rect -192 -145 -124 -111
rect -34 -145 34 -111
rect 124 -145 192 -111
rect 282 -145 350 -111
rect 440 -145 508 -111
rect 598 -145 666 -111
rect 756 -145 824 -111
rect 914 -145 982 -111
<< locali >>
rect -1158 214 -1062 248
rect 1062 214 1158 248
rect -1158 151 -1124 214
rect 1124 151 1158 214
rect -1044 124 -1010 140
rect -1044 -68 -1010 -52
rect -886 124 -852 140
rect -886 -68 -852 -52
rect -728 124 -694 140
rect -728 -68 -694 -52
rect -570 124 -536 140
rect -570 -68 -536 -52
rect -412 124 -378 140
rect -412 -68 -378 -52
rect -254 124 -220 140
rect -254 -68 -220 -52
rect -96 124 -62 140
rect -96 -68 -62 -52
rect 62 124 96 140
rect 62 -68 96 -52
rect 220 124 254 140
rect 220 -68 254 -52
rect 378 124 412 140
rect 378 -68 412 -52
rect 536 124 570 140
rect 536 -68 570 -52
rect 694 124 728 140
rect 694 -68 728 -52
rect 852 124 886 140
rect 852 -68 886 -52
rect 1010 124 1044 140
rect 1010 -68 1044 -52
rect -998 -145 -982 -111
rect -914 -145 -898 -111
rect -840 -145 -824 -111
rect -756 -145 -740 -111
rect -682 -145 -666 -111
rect -598 -145 -582 -111
rect -524 -145 -508 -111
rect -440 -145 -424 -111
rect -366 -145 -350 -111
rect -282 -145 -266 -111
rect -208 -145 -192 -111
rect -124 -145 -108 -111
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect 108 -145 124 -111
rect 192 -145 208 -111
rect 266 -145 282 -111
rect 350 -145 366 -111
rect 424 -145 440 -111
rect 508 -145 524 -111
rect 582 -145 598 -111
rect 666 -145 682 -111
rect 740 -145 756 -111
rect 824 -145 840 -111
rect 898 -145 914 -111
rect 982 -145 998 -111
rect -1158 -214 -1124 -151
rect 1124 -214 1158 -151
rect -1158 -248 -1062 -214
rect 1062 -248 1158 -214
<< viali >>
rect -1044 -52 -1010 124
rect -886 -52 -852 124
rect -728 -52 -694 124
rect -570 -52 -536 124
rect -412 -52 -378 124
rect -254 -52 -220 124
rect -96 -52 -62 124
rect 62 -52 96 124
rect 220 -52 254 124
rect 378 -52 412 124
rect 536 -52 570 124
rect 694 -52 728 124
rect 852 -52 886 124
rect 1010 -52 1044 124
rect -982 -145 -914 -111
rect -824 -145 -756 -111
rect -666 -145 -598 -111
rect -508 -145 -440 -111
rect -350 -145 -282 -111
rect -192 -145 -124 -111
rect -34 -145 34 -111
rect 124 -145 192 -111
rect 282 -145 350 -111
rect 440 -145 508 -111
rect 598 -145 666 -111
rect 756 -145 824 -111
rect 914 -145 982 -111
<< metal1 >>
rect -1050 124 -1004 136
rect -1050 -52 -1044 124
rect -1010 -52 -1004 124
rect -1050 -64 -1004 -52
rect -892 124 -846 136
rect -892 -52 -886 124
rect -852 -52 -846 124
rect -892 -64 -846 -52
rect -734 124 -688 136
rect -734 -52 -728 124
rect -694 -52 -688 124
rect -734 -64 -688 -52
rect -576 124 -530 136
rect -576 -52 -570 124
rect -536 -52 -530 124
rect -576 -64 -530 -52
rect -418 124 -372 136
rect -418 -52 -412 124
rect -378 -52 -372 124
rect -418 -64 -372 -52
rect -260 124 -214 136
rect -260 -52 -254 124
rect -220 -52 -214 124
rect -260 -64 -214 -52
rect -102 124 -56 136
rect -102 -52 -96 124
rect -62 -52 -56 124
rect -102 -64 -56 -52
rect 56 124 102 136
rect 56 -52 62 124
rect 96 -52 102 124
rect 56 -64 102 -52
rect 214 124 260 136
rect 214 -52 220 124
rect 254 -52 260 124
rect 214 -64 260 -52
rect 372 124 418 136
rect 372 -52 378 124
rect 412 -52 418 124
rect 372 -64 418 -52
rect 530 124 576 136
rect 530 -52 536 124
rect 570 -52 576 124
rect 530 -64 576 -52
rect 688 124 734 136
rect 688 -52 694 124
rect 728 -52 734 124
rect 688 -64 734 -52
rect 846 124 892 136
rect 846 -52 852 124
rect 886 -52 892 124
rect 846 -64 892 -52
rect 1004 124 1050 136
rect 1004 -52 1010 124
rect 1044 -52 1050 124
rect 1004 -64 1050 -52
rect -994 -111 -902 -105
rect -994 -145 -982 -111
rect -914 -145 -902 -111
rect -994 -151 -902 -145
rect -836 -111 -744 -105
rect -836 -145 -824 -111
rect -756 -145 -744 -111
rect -836 -151 -744 -145
rect -678 -111 -586 -105
rect -678 -145 -666 -111
rect -598 -145 -586 -111
rect -678 -151 -586 -145
rect -520 -111 -428 -105
rect -520 -145 -508 -111
rect -440 -145 -428 -111
rect -520 -151 -428 -145
rect -362 -111 -270 -105
rect -362 -145 -350 -111
rect -282 -145 -270 -111
rect -362 -151 -270 -145
rect -204 -111 -112 -105
rect -204 -145 -192 -111
rect -124 -145 -112 -111
rect -204 -151 -112 -145
rect -46 -111 46 -105
rect -46 -145 -34 -111
rect 34 -145 46 -111
rect -46 -151 46 -145
rect 112 -111 204 -105
rect 112 -145 124 -111
rect 192 -145 204 -111
rect 112 -151 204 -145
rect 270 -111 362 -105
rect 270 -145 282 -111
rect 350 -145 362 -111
rect 270 -151 362 -145
rect 428 -111 520 -105
rect 428 -145 440 -111
rect 508 -145 520 -111
rect 428 -151 520 -145
rect 586 -111 678 -105
rect 586 -145 598 -111
rect 666 -145 678 -111
rect 586 -151 678 -145
rect 744 -111 836 -105
rect 744 -145 756 -111
rect 824 -145 836 -111
rect 744 -151 836 -145
rect 902 -111 994 -105
rect 902 -145 914 -111
rect 982 -145 994 -111
rect 902 -151 994 -145
<< properties >>
string FIXED_BBOX -1141 -231 1141 231
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

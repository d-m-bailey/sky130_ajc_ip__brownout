magic
tech sky130A
magscale 1 2
timestamp 1712784588
<< nwell >>
rect -154 -198 154 164
<< pmos >>
rect -60 -136 60 64
<< pdiff >>
rect -118 52 -60 64
rect -118 -124 -106 52
rect -72 -124 -60 52
rect -118 -136 -60 -124
rect 60 52 118 64
rect 60 -124 72 52
rect 106 -124 118 52
rect 60 -136 118 -124
<< pdiffc >>
rect -106 -124 -72 52
rect 72 -124 106 52
<< poly >>
rect -60 145 60 161
rect -60 111 -44 145
rect 44 111 60 145
rect -60 64 60 111
rect -60 -162 60 -136
<< polycont >>
rect -44 111 44 145
<< locali >>
rect -60 111 -44 145
rect 44 111 60 145
rect -106 52 -72 68
rect -106 -140 -72 -124
rect 72 52 106 68
rect 72 -140 106 -124
<< viali >>
rect -44 111 44 145
rect -106 -124 -72 52
rect 72 -124 106 52
<< metal1 >>
rect -56 145 56 151
rect -56 111 -44 145
rect 44 111 56 145
rect -56 105 56 111
rect -112 52 -66 64
rect -112 -124 -106 52
rect -72 -124 -66 52
rect -112 -136 -66 -124
rect 66 52 112 64
rect 66 -124 72 52
rect 106 -124 112 52
rect 66 -136 112 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

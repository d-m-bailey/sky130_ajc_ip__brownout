** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__brownout/cace/trip_up_down.sch
**.subckt trip_up_down
Ibias vbp GND 200n
XM1 ibg_200n vbp avdd_bg avdd_bg sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM0 vbp vbp avdd_bg avdd_bg sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 itest GND 1e6 m=1
C1 outb GND 20p m=1
xIbrout avdd avss outb dvdd osc_ck dvss dcomp vbg_1v2 otrip[2] otrip[1] otrip[0] itest brout_filt vtrip[2] vtrip[1] vtrip[0]  vin_brout ena force_ena_rc_osc vin_vunder force_dis_rc_osc timed_out vunder force_short_oneshot isrc_sel ibg_200n sky130_ajc_ip__brownout
Vavss avss GND DC 0
Vena ena GND DC 1.8
Vavdd avdd GND pwl (0 2 3m 3.6 6m 2) DC 3.3
.save i(vavdd)
Vbg1v2 vbg_1v2 GND DC 1.2
Vdvss dvss GND DC 0
Vdvdd dvdd GND DC 1.8
.save i(vdvdd)
Vvotrip0 otrip[0] GND DC 0.0
.save i(vvotrip0)
Vvotrip1 otrip[1] GND DC 0.0
.save i(vvotrip1)
Vvotrip2 otrip[2] GND DC 1.8
.save i(vvotrip2)
Vvotrip3 otrip[3] GND DC 0.0
.save i(vvotrip3)
Visrc_sel isrc_sel GND DC 0.0
Vvvtrip0 vtrip[0] GND DC 0.0
.save i(vvvtrip0)
Vvvtrip1 vtrip[1] GND DC 0.0
.save i(vvvtrip1)
Vvvtrip2 vtrip[2] GND DC 1.8
.save i(vvvtrip2)
Vvvtrip3 vtrip[3] GND DC 0.0
.save i(vvvtrip3)
Vforce_dis_rc_osc force_dis_rc_osc GND DC 1.8
Vforce_short_oneshot force_short_oneshot GND DC 0.0
Vavdd_bg avdd_bg GND DC 3.3
Vforce_ena_rc_osc force_ena_rc_osc GND DC 0.0
**** begin user architecture code

* CACE gensim simulation file hysteresis_br_8
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find trip voltage by ramping Vavdd, both up and down.

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
*.include ./netlist/schematic/sky130_ajc_ip__brownout.spice


.option TEMP=85
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
*.option reltol=5e-5
.option reltol=1e-3
.option abstol=1e-3

.save all



.csparam dvdd2=0.9
.control
tran 1u 6m
meas tran otrip_r find v(avdd) when v(dcomp)=$&dvdd2 td=3m rise=1
meas tran otrip_f find v(avdd) when v(dcomp)=$&dvdd2 td=300u fall=1
meas tran vtrip_r find v(avdd) when v(vunder)=$&dvdd2 td=300u rise=1
meas tran vtrip_f find v(avdd) when v(vunder)=$&dvdd2 td=3m fall=1
echo $&otrip_r > ngspice/hysteresis_br_8.data
echo $&otrip_f >> ngspice/hysteresis_br_8.data
echo $&vtrip_r >> ngspice/hysteresis_br_8.data
echo $&vtrip_f >> ngspice/hysteresis_br_8.data
quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  xschem/sky130_ajc_ip__brownout.sym # of pins=22
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__brownout/xschem/sky130_ajc_ip__brownout.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__brownout/xschem/sky130_ajc_ip__brownout.sch
.subckt sky130_ajc_ip__brownout avdd avss outb dvdd osc_ck dvss dcomp vbg_1v2 otrip[2] otrip[1] otrip[0] itest brout_filt vtrip[2] vtrip[1] vtrip[0] vin_brout ena force_ena_rc_osc vin_vunder force_dis_rc_osc timed_out vunder force_short_oneshot isrc_sel ibg_200n
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin vbg_1v2
*.ipin otrip[2],otrip[1],otrip[0]
*.ipin ena
*.ipin force_dis_rc_osc
*.ipin force_short_oneshot
*.ipin isrc_sel
*.ipin ibg_200n
*.opin vin_brout
*.opin outb
*.opin osc_ck
*.opin brout_filt
*.opin itest
*.opin timed_out
*.ipin vtrip[2],vtrip[1],vtrip[0]
*.opin vin_vunder
*.opin vunder
*.ipin force_ena_rc_osc
*.opin dcomp
xIana vin_brout otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_ otrip_decoded_1_ otrip_decoded_0_ vin_vunder vbg_1v2 ena avdd ibg_200n itest avss dvdd isrc_sel dvss vtrip_decoded_7_ vtrip_decoded_6_ vtrip_decoded_5_ vtrip_decoded_4_ vtrip_decoded_3_ vtrip_decoded_2_ vtrip_decoded_1_ vtrip_decoded_0_ dcomp brout_filt osc_ck osc_ena vunder outb outb_unbuf brownout_ana_rcx
**** begin user architecture code



r0 otrip[0] otrip0 1
r1 otrip[1] otrip1 1
r2 otrip[2] otrip2 1
r3 vtrip[0] vtrip0 1
r4 vtrip[1] vtrip1 1
r5 vtrip[2] vtrip2 1

*XSPICE CO-SIM netlist
.include brownout_dig.out.spice
xibrownout_dig dvss dvdd brout_filt dcomp ena force_dis_rc_osc force_ena_rc_osc force_short_oneshot osc_ck osc_ena otrip0 otrip1 otrip2 otrip_decoded_0_ otrip_decoded_1_ otrip_decoded_2_ otrip_decoded_3_ otrip_decoded_4_ otrip_decoded_5_ otrip_decoded_6_ otrip_decoded_7_ outb_unbuf timed_out vtrip0 vtrip1 vtrip2 vtrip_decoded_0_ vtrip_decoded_1_ vtrip_decoded_2_ vtrip_decoded_3_ vtrip_decoded_4_ vtrip_decoded_5_ vtrip_decoded_6_ vtrip_decoded_7_ brownout_dig


**** end user architecture code
.ends


* expanding   symbol:  xschem/brownout_ana_rcx.sym # of pins=20
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__brownout/xschem/brownout_ana_rcx.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__brownout/xschem/brownout_ana_rcx.sch
.subckt brownout_ana_rcx vin_brout otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3] otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vin_vunder vbg_1v2 ena avdd ibg_200n itest avss dvdd isrc_sel dvss vtrip_decoded[7] vtrip_decoded[6] vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2] vtrip_decoded[1] vtrip_decoded[0] dcomp brout_filt osc_ck osc_ena vunder outb outb_unbuf
*.ipin vbg_1v2
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin ena
*.ipin isrc_sel
*.ipin ibg_200n
*.opin dcomp
*.opin itest
*.ipin osc_ena
*.opin osc_ck
*.ipin otrip_decoded[7],otrip_decoded[6],otrip_decoded[5],otrip_decoded[4],otrip_decoded[3],otrip_decoded[2],otrip_decoded[1],otrip_decoded[0]
*.opin vin_brout
*.ipin outb_unbuf
*.opin outb
*.opin vunder
*.ipin vtrip_decoded[7],vtrip_decoded[6],vtrip_decoded[5],vtrip_decoded[4],vtrip_decoded[3],vtrip_decoded[2],vtrip_decoded[1],vtrip_decoded[0]
*.opin vin_vunder
*.opin brout_filt
**** begin user architecture code



.include mag/rcx/brownout_ana_rcx.spice

xIana vin_brout otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3] otrip_decoded[2]  otrip_decoded[1] otrip_decoded[0] vin_vunder vbg_1v2 ena avdd ibg_200n itest avss dvdd isrc_sel dvss vtrip_decoded[7] vtrip_decoded[6]  vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2] vtrip_decoded[1] vtrip_decoded[0] dcomp brout_filt osc_ck osc_ena vunder outb  outb_unbuf brownout_ana



**** end user architecture code
.ends

.GLOBAL GND
.end

magic
tech sky130A
magscale 1 2
timestamp 1712722749
<< nwell >>
rect -1194 -319 1194 319
<< pmos >>
rect -998 -100 -898 100
rect -840 -100 -740 100
rect -682 -100 -582 100
rect -524 -100 -424 100
rect -366 -100 -266 100
rect -208 -100 -108 100
rect -50 -100 50 100
rect 108 -100 208 100
rect 266 -100 366 100
rect 424 -100 524 100
rect 582 -100 682 100
rect 740 -100 840 100
rect 898 -100 998 100
<< pdiff >>
rect -1056 88 -998 100
rect -1056 -88 -1044 88
rect -1010 -88 -998 88
rect -1056 -100 -998 -88
rect -898 88 -840 100
rect -898 -88 -886 88
rect -852 -88 -840 88
rect -898 -100 -840 -88
rect -740 88 -682 100
rect -740 -88 -728 88
rect -694 -88 -682 88
rect -740 -100 -682 -88
rect -582 88 -524 100
rect -582 -88 -570 88
rect -536 -88 -524 88
rect -582 -100 -524 -88
rect -424 88 -366 100
rect -424 -88 -412 88
rect -378 -88 -366 88
rect -424 -100 -366 -88
rect -266 88 -208 100
rect -266 -88 -254 88
rect -220 -88 -208 88
rect -266 -100 -208 -88
rect -108 88 -50 100
rect -108 -88 -96 88
rect -62 -88 -50 88
rect -108 -100 -50 -88
rect 50 88 108 100
rect 50 -88 62 88
rect 96 -88 108 88
rect 50 -100 108 -88
rect 208 88 266 100
rect 208 -88 220 88
rect 254 -88 266 88
rect 208 -100 266 -88
rect 366 88 424 100
rect 366 -88 378 88
rect 412 -88 424 88
rect 366 -100 424 -88
rect 524 88 582 100
rect 524 -88 536 88
rect 570 -88 582 88
rect 524 -100 582 -88
rect 682 88 740 100
rect 682 -88 694 88
rect 728 -88 740 88
rect 682 -100 740 -88
rect 840 88 898 100
rect 840 -88 852 88
rect 886 -88 898 88
rect 840 -100 898 -88
rect 998 88 1056 100
rect 998 -88 1010 88
rect 1044 -88 1056 88
rect 998 -100 1056 -88
<< pdiffc >>
rect -1044 -88 -1010 88
rect -886 -88 -852 88
rect -728 -88 -694 88
rect -570 -88 -536 88
rect -412 -88 -378 88
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
rect 378 -88 412 88
rect 536 -88 570 88
rect 694 -88 728 88
rect 852 -88 886 88
rect 1010 -88 1044 88
<< nsubdiff >>
rect -1158 249 -1062 283
rect 1062 249 1158 283
rect -1158 187 -1124 249
rect 1124 187 1158 249
rect -1158 -249 -1124 -187
rect 1124 -249 1158 -187
rect -1158 -283 -1062 -249
rect 1062 -283 1158 -249
<< nsubdiffcont >>
rect -1062 249 1062 283
rect -1158 -187 -1124 187
rect 1124 -187 1158 187
rect -1062 -283 1062 -249
<< poly >>
rect -998 181 -898 197
rect -998 147 -982 181
rect -914 147 -898 181
rect -998 100 -898 147
rect -840 181 -740 197
rect -840 147 -824 181
rect -756 147 -740 181
rect -840 100 -740 147
rect -682 181 -582 197
rect -682 147 -666 181
rect -598 147 -582 181
rect -682 100 -582 147
rect -524 181 -424 197
rect -524 147 -508 181
rect -440 147 -424 181
rect -524 100 -424 147
rect -366 181 -266 197
rect -366 147 -350 181
rect -282 147 -266 181
rect -366 100 -266 147
rect -208 181 -108 197
rect -208 147 -192 181
rect -124 147 -108 181
rect -208 100 -108 147
rect -50 181 50 197
rect -50 147 -34 181
rect 34 147 50 181
rect -50 100 50 147
rect 108 181 208 197
rect 108 147 124 181
rect 192 147 208 181
rect 108 100 208 147
rect 266 181 366 197
rect 266 147 282 181
rect 350 147 366 181
rect 266 100 366 147
rect 424 181 524 197
rect 424 147 440 181
rect 508 147 524 181
rect 424 100 524 147
rect 582 181 682 197
rect 582 147 598 181
rect 666 147 682 181
rect 582 100 682 147
rect 740 181 840 197
rect 740 147 756 181
rect 824 147 840 181
rect 740 100 840 147
rect 898 181 998 197
rect 898 147 914 181
rect 982 147 998 181
rect 898 100 998 147
rect -998 -147 -898 -100
rect -998 -181 -982 -147
rect -914 -181 -898 -147
rect -998 -197 -898 -181
rect -840 -147 -740 -100
rect -840 -181 -824 -147
rect -756 -181 -740 -147
rect -840 -197 -740 -181
rect -682 -147 -582 -100
rect -682 -181 -666 -147
rect -598 -181 -582 -147
rect -682 -197 -582 -181
rect -524 -147 -424 -100
rect -524 -181 -508 -147
rect -440 -181 -424 -147
rect -524 -197 -424 -181
rect -366 -147 -266 -100
rect -366 -181 -350 -147
rect -282 -181 -266 -147
rect -366 -197 -266 -181
rect -208 -147 -108 -100
rect -208 -181 -192 -147
rect -124 -181 -108 -147
rect -208 -197 -108 -181
rect -50 -147 50 -100
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect -50 -197 50 -181
rect 108 -147 208 -100
rect 108 -181 124 -147
rect 192 -181 208 -147
rect 108 -197 208 -181
rect 266 -147 366 -100
rect 266 -181 282 -147
rect 350 -181 366 -147
rect 266 -197 366 -181
rect 424 -147 524 -100
rect 424 -181 440 -147
rect 508 -181 524 -147
rect 424 -197 524 -181
rect 582 -147 682 -100
rect 582 -181 598 -147
rect 666 -181 682 -147
rect 582 -197 682 -181
rect 740 -147 840 -100
rect 740 -181 756 -147
rect 824 -181 840 -147
rect 740 -197 840 -181
rect 898 -147 998 -100
rect 898 -181 914 -147
rect 982 -181 998 -147
rect 898 -197 998 -181
<< polycont >>
rect -982 147 -914 181
rect -824 147 -756 181
rect -666 147 -598 181
rect -508 147 -440 181
rect -350 147 -282 181
rect -192 147 -124 181
rect -34 147 34 181
rect 124 147 192 181
rect 282 147 350 181
rect 440 147 508 181
rect 598 147 666 181
rect 756 147 824 181
rect 914 147 982 181
rect -982 -181 -914 -147
rect -824 -181 -756 -147
rect -666 -181 -598 -147
rect -508 -181 -440 -147
rect -350 -181 -282 -147
rect -192 -181 -124 -147
rect -34 -181 34 -147
rect 124 -181 192 -147
rect 282 -181 350 -147
rect 440 -181 508 -147
rect 598 -181 666 -147
rect 756 -181 824 -147
rect 914 -181 982 -147
<< locali >>
rect -1158 249 -1062 283
rect 1062 249 1158 283
rect -1158 187 -1124 249
rect 1124 187 1158 249
rect -998 147 -982 181
rect -914 147 -898 181
rect -840 147 -824 181
rect -756 147 -740 181
rect -682 147 -666 181
rect -598 147 -582 181
rect -524 147 -508 181
rect -440 147 -424 181
rect -366 147 -350 181
rect -282 147 -266 181
rect -208 147 -192 181
rect -124 147 -108 181
rect -50 147 -34 181
rect 34 147 50 181
rect 108 147 124 181
rect 192 147 208 181
rect 266 147 282 181
rect 350 147 366 181
rect 424 147 440 181
rect 508 147 524 181
rect 582 147 598 181
rect 666 147 682 181
rect 740 147 756 181
rect 824 147 840 181
rect 898 147 914 181
rect 982 147 998 181
rect -1044 88 -1010 104
rect -1044 -104 -1010 -88
rect -886 88 -852 104
rect -886 -104 -852 -88
rect -728 88 -694 104
rect -728 -104 -694 -88
rect -570 88 -536 104
rect -570 -104 -536 -88
rect -412 88 -378 104
rect -412 -104 -378 -88
rect -254 88 -220 104
rect -254 -104 -220 -88
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect 220 88 254 104
rect 220 -104 254 -88
rect 378 88 412 104
rect 378 -104 412 -88
rect 536 88 570 104
rect 536 -104 570 -88
rect 694 88 728 104
rect 694 -104 728 -88
rect 852 88 886 104
rect 852 -104 886 -88
rect 1010 88 1044 104
rect 1010 -104 1044 -88
rect -998 -181 -982 -147
rect -914 -181 -898 -147
rect -840 -181 -824 -147
rect -756 -181 -740 -147
rect -682 -181 -666 -147
rect -598 -181 -582 -147
rect -524 -181 -508 -147
rect -440 -181 -424 -147
rect -366 -181 -350 -147
rect -282 -181 -266 -147
rect -208 -181 -192 -147
rect -124 -181 -108 -147
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect 108 -181 124 -147
rect 192 -181 208 -147
rect 266 -181 282 -147
rect 350 -181 366 -147
rect 424 -181 440 -147
rect 508 -181 524 -147
rect 582 -181 598 -147
rect 666 -181 682 -147
rect 740 -181 756 -147
rect 824 -181 840 -147
rect 898 -181 914 -147
rect 982 -181 998 -147
rect -1158 -249 -1124 -187
rect 1124 -249 1158 -187
rect -1158 -283 -1062 -249
rect 1062 -283 1158 -249
<< viali >>
rect -982 147 -914 181
rect -824 147 -756 181
rect -666 147 -598 181
rect -508 147 -440 181
rect -350 147 -282 181
rect -192 147 -124 181
rect -34 147 34 181
rect 124 147 192 181
rect 282 147 350 181
rect 440 147 508 181
rect 598 147 666 181
rect 756 147 824 181
rect 914 147 982 181
rect -1044 -88 -1010 88
rect -886 -88 -852 88
rect -728 -88 -694 88
rect -570 -88 -536 88
rect -412 -88 -378 88
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
rect 378 -88 412 88
rect 536 -88 570 88
rect 694 -88 728 88
rect 852 -88 886 88
rect 1010 -88 1044 88
rect -982 -181 -914 -147
rect -824 -181 -756 -147
rect -666 -181 -598 -147
rect -508 -181 -440 -147
rect -350 -181 -282 -147
rect -192 -181 -124 -147
rect -34 -181 34 -147
rect 124 -181 192 -147
rect 282 -181 350 -147
rect 440 -181 508 -147
rect 598 -181 666 -147
rect 756 -181 824 -147
rect 914 -181 982 -147
<< metal1 >>
rect -994 181 -902 187
rect -994 147 -982 181
rect -914 147 -902 181
rect -994 141 -902 147
rect -836 181 -744 187
rect -836 147 -824 181
rect -756 147 -744 181
rect -836 141 -744 147
rect -678 181 -586 187
rect -678 147 -666 181
rect -598 147 -586 181
rect -678 141 -586 147
rect -520 181 -428 187
rect -520 147 -508 181
rect -440 147 -428 181
rect -520 141 -428 147
rect -362 181 -270 187
rect -362 147 -350 181
rect -282 147 -270 181
rect -362 141 -270 147
rect -204 181 -112 187
rect -204 147 -192 181
rect -124 147 -112 181
rect -204 141 -112 147
rect -46 181 46 187
rect -46 147 -34 181
rect 34 147 46 181
rect -46 141 46 147
rect 112 181 204 187
rect 112 147 124 181
rect 192 147 204 181
rect 112 141 204 147
rect 270 181 362 187
rect 270 147 282 181
rect 350 147 362 181
rect 270 141 362 147
rect 428 181 520 187
rect 428 147 440 181
rect 508 147 520 181
rect 428 141 520 147
rect 586 181 678 187
rect 586 147 598 181
rect 666 147 678 181
rect 586 141 678 147
rect 744 181 836 187
rect 744 147 756 181
rect 824 147 836 181
rect 744 141 836 147
rect 902 181 994 187
rect 902 147 914 181
rect 982 147 994 181
rect 902 141 994 147
rect -1050 88 -1004 100
rect -1050 -88 -1044 88
rect -1010 -88 -1004 88
rect -1050 -100 -1004 -88
rect -892 88 -846 100
rect -892 -88 -886 88
rect -852 -88 -846 88
rect -892 -100 -846 -88
rect -734 88 -688 100
rect -734 -88 -728 88
rect -694 -88 -688 88
rect -734 -100 -688 -88
rect -576 88 -530 100
rect -576 -88 -570 88
rect -536 -88 -530 88
rect -576 -100 -530 -88
rect -418 88 -372 100
rect -418 -88 -412 88
rect -378 -88 -372 88
rect -418 -100 -372 -88
rect -260 88 -214 100
rect -260 -88 -254 88
rect -220 -88 -214 88
rect -260 -100 -214 -88
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect 214 88 260 100
rect 214 -88 220 88
rect 254 -88 260 88
rect 214 -100 260 -88
rect 372 88 418 100
rect 372 -88 378 88
rect 412 -88 418 88
rect 372 -100 418 -88
rect 530 88 576 100
rect 530 -88 536 88
rect 570 -88 576 88
rect 530 -100 576 -88
rect 688 88 734 100
rect 688 -88 694 88
rect 728 -88 734 88
rect 688 -100 734 -88
rect 846 88 892 100
rect 846 -88 852 88
rect 886 -88 892 88
rect 846 -100 892 -88
rect 1004 88 1050 100
rect 1004 -88 1010 88
rect 1044 -88 1050 88
rect 1004 -100 1050 -88
rect -994 -147 -902 -141
rect -994 -181 -982 -147
rect -914 -181 -902 -147
rect -994 -187 -902 -181
rect -836 -147 -744 -141
rect -836 -181 -824 -147
rect -756 -181 -744 -147
rect -836 -187 -744 -181
rect -678 -147 -586 -141
rect -678 -181 -666 -147
rect -598 -181 -586 -147
rect -678 -187 -586 -181
rect -520 -147 -428 -141
rect -520 -181 -508 -147
rect -440 -181 -428 -147
rect -520 -187 -428 -181
rect -362 -147 -270 -141
rect -362 -181 -350 -147
rect -282 -181 -270 -147
rect -362 -187 -270 -181
rect -204 -147 -112 -141
rect -204 -181 -192 -147
rect -124 -181 -112 -147
rect -204 -187 -112 -181
rect -46 -147 46 -141
rect -46 -181 -34 -147
rect 34 -181 46 -147
rect -46 -187 46 -181
rect 112 -147 204 -141
rect 112 -181 124 -147
rect 192 -181 204 -147
rect 112 -187 204 -181
rect 270 -147 362 -141
rect 270 -181 282 -147
rect 350 -181 362 -147
rect 270 -187 362 -181
rect 428 -147 520 -141
rect 428 -181 440 -147
rect 508 -181 520 -147
rect 428 -187 520 -181
rect 586 -147 678 -141
rect 586 -181 598 -147
rect 666 -181 678 -147
rect 586 -187 678 -181
rect 744 -147 836 -141
rect 744 -181 756 -147
rect 824 -181 836 -147
rect 744 -187 836 -181
rect 902 -147 994 -141
rect 902 -181 914 -147
rect 982 -181 994 -147
rect 902 -187 994 -181
<< properties >>
string FIXED_BBOX -1141 -266 1141 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712722749
<< nwell >>
rect -539 -164 539 198
<< pmos >>
rect -445 -64 -345 136
rect -287 -64 -187 136
rect -129 -64 -29 136
rect 29 -64 129 136
rect 187 -64 287 136
rect 345 -64 445 136
<< pdiff >>
rect -503 124 -445 136
rect -503 -52 -491 124
rect -457 -52 -445 124
rect -503 -64 -445 -52
rect -345 124 -287 136
rect -345 -52 -333 124
rect -299 -52 -287 124
rect -345 -64 -287 -52
rect -187 124 -129 136
rect -187 -52 -175 124
rect -141 -52 -129 124
rect -187 -64 -129 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 129 124 187 136
rect 129 -52 141 124
rect 175 -52 187 124
rect 129 -64 187 -52
rect 287 124 345 136
rect 287 -52 299 124
rect 333 -52 345 124
rect 287 -64 345 -52
rect 445 124 503 136
rect 445 -52 457 124
rect 491 -52 503 124
rect 445 -64 503 -52
<< pdiffc >>
rect -491 -52 -457 124
rect -333 -52 -299 124
rect -175 -52 -141 124
rect -17 -52 17 124
rect 141 -52 175 124
rect 299 -52 333 124
rect 457 -52 491 124
<< poly >>
rect -445 136 -345 162
rect -287 136 -187 162
rect -129 136 -29 162
rect 29 136 129 162
rect 187 136 287 162
rect 345 136 445 162
rect -445 -111 -345 -64
rect -445 -145 -429 -111
rect -361 -145 -345 -111
rect -445 -161 -345 -145
rect -287 -111 -187 -64
rect -287 -145 -271 -111
rect -203 -145 -187 -111
rect -287 -161 -187 -145
rect -129 -111 -29 -64
rect -129 -145 -113 -111
rect -45 -145 -29 -111
rect -129 -161 -29 -145
rect 29 -111 129 -64
rect 29 -145 45 -111
rect 113 -145 129 -111
rect 29 -161 129 -145
rect 187 -111 287 -64
rect 187 -145 203 -111
rect 271 -145 287 -111
rect 187 -161 287 -145
rect 345 -111 445 -64
rect 345 -145 361 -111
rect 429 -145 445 -111
rect 345 -161 445 -145
<< polycont >>
rect -429 -145 -361 -111
rect -271 -145 -203 -111
rect -113 -145 -45 -111
rect 45 -145 113 -111
rect 203 -145 271 -111
rect 361 -145 429 -111
<< locali >>
rect -491 124 -457 140
rect -491 -68 -457 -52
rect -333 124 -299 140
rect -333 -68 -299 -52
rect -175 124 -141 140
rect -175 -68 -141 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 141 124 175 140
rect 141 -68 175 -52
rect 299 124 333 140
rect 299 -68 333 -52
rect 457 124 491 140
rect 457 -68 491 -52
rect -445 -145 -429 -111
rect -361 -145 -345 -111
rect -287 -145 -271 -111
rect -203 -145 -187 -111
rect -129 -145 -113 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 113 -145 129 -111
rect 187 -145 203 -111
rect 271 -145 287 -111
rect 345 -145 361 -111
rect 429 -145 445 -111
<< viali >>
rect -491 -52 -457 124
rect -333 -52 -299 124
rect -175 -52 -141 124
rect -17 -52 17 124
rect 141 -52 175 124
rect 299 -52 333 124
rect 457 -52 491 124
rect -429 -145 -361 -111
rect -271 -145 -203 -111
rect -113 -145 -45 -111
rect 45 -145 113 -111
rect 203 -145 271 -111
rect 361 -145 429 -111
<< metal1 >>
rect -497 124 -451 136
rect -497 -52 -491 124
rect -457 -52 -451 124
rect -497 -64 -451 -52
rect -339 124 -293 136
rect -339 -52 -333 124
rect -299 -52 -293 124
rect -339 -64 -293 -52
rect -181 124 -135 136
rect -181 -52 -175 124
rect -141 -52 -135 124
rect -181 -64 -135 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 135 124 181 136
rect 135 -52 141 124
rect 175 -52 181 124
rect 135 -64 181 -52
rect 293 124 339 136
rect 293 -52 299 124
rect 333 -52 339 124
rect 293 -64 339 -52
rect 451 124 497 136
rect 451 -52 457 124
rect 491 -52 497 124
rect 451 -64 497 -52
rect -441 -111 -349 -105
rect -441 -145 -429 -111
rect -361 -145 -349 -111
rect -441 -151 -349 -145
rect -283 -111 -191 -105
rect -283 -145 -271 -111
rect -203 -145 -191 -111
rect -283 -151 -191 -145
rect -125 -111 -33 -105
rect -125 -145 -113 -111
rect -45 -145 -33 -111
rect -125 -151 -33 -145
rect 33 -111 125 -105
rect 33 -145 45 -111
rect 113 -145 125 -111
rect 33 -151 125 -145
rect 191 -111 283 -105
rect 191 -145 203 -111
rect 271 -145 283 -111
rect 191 -151 283 -145
rect 349 -111 441 -105
rect 349 -145 361 -111
rect 429 -145 441 -111
rect 349 -151 441 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

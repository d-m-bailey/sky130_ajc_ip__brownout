magic
tech sky130A
magscale 1 2
timestamp 1712722749
<< nmos >>
rect -287 -131 -187 69
rect -129 -131 -29 69
rect 29 -131 129 69
rect 187 -131 287 69
<< ndiff >>
rect -345 57 -287 69
rect -345 -119 -333 57
rect -299 -119 -287 57
rect -345 -131 -287 -119
rect -187 57 -129 69
rect -187 -119 -175 57
rect -141 -119 -129 57
rect -187 -131 -129 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 129 57 187 69
rect 129 -119 141 57
rect 175 -119 187 57
rect 129 -131 187 -119
rect 287 57 345 69
rect 287 -119 299 57
rect 333 -119 345 57
rect 287 -131 345 -119
<< ndiffc >>
rect -333 -119 -299 57
rect -175 -119 -141 57
rect -17 -119 17 57
rect 141 -119 175 57
rect 299 -119 333 57
<< poly >>
rect -287 141 -187 157
rect -287 107 -271 141
rect -203 107 -187 141
rect -287 69 -187 107
rect -129 141 -29 157
rect -129 107 -113 141
rect -45 107 -29 141
rect -129 69 -29 107
rect 29 141 129 157
rect 29 107 45 141
rect 113 107 129 141
rect 29 69 129 107
rect 187 141 287 157
rect 187 107 203 141
rect 271 107 287 141
rect 187 69 287 107
rect -287 -157 -187 -131
rect -129 -157 -29 -131
rect 29 -157 129 -131
rect 187 -157 287 -131
<< polycont >>
rect -271 107 -203 141
rect -113 107 -45 141
rect 45 107 113 141
rect 203 107 271 141
<< locali >>
rect -287 107 -271 141
rect -203 107 -187 141
rect -129 107 -113 141
rect -45 107 -29 141
rect 29 107 45 141
rect 113 107 129 141
rect 187 107 203 141
rect 271 107 287 141
rect -333 57 -299 73
rect -333 -135 -299 -119
rect -175 57 -141 73
rect -175 -135 -141 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 141 57 175 73
rect 141 -135 175 -119
rect 299 57 333 73
rect 299 -135 333 -119
<< viali >>
rect -271 107 -203 141
rect -113 107 -45 141
rect 45 107 113 141
rect 203 107 271 141
rect -333 -119 -299 57
rect -175 -119 -141 57
rect -17 -119 17 57
rect 141 -119 175 57
rect 299 -119 333 57
<< metal1 >>
rect -283 141 -191 147
rect -283 107 -271 141
rect -203 107 -191 141
rect -283 101 -191 107
rect -125 141 -33 147
rect -125 107 -113 141
rect -45 107 -33 141
rect -125 101 -33 107
rect 33 141 125 147
rect 33 107 45 141
rect 113 107 125 141
rect 33 101 125 107
rect 191 141 283 147
rect 191 107 203 141
rect 271 107 283 141
rect 191 101 283 107
rect -339 57 -293 69
rect -339 -119 -333 57
rect -299 -119 -293 57
rect -339 -131 -293 -119
rect -181 57 -135 69
rect -181 -119 -175 57
rect -141 -119 -135 57
rect -181 -131 -135 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 135 57 181 69
rect 135 -119 141 57
rect 175 -119 181 57
rect 135 -131 181 -119
rect 293 57 339 69
rect 293 -119 299 57
rect 333 -119 339 57
rect 293 -131 339 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

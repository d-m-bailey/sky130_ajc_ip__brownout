magic
tech sky130A
magscale 1 2
timestamp 1712930986
<< nwell >>
rect -358 -909 358 909
<< mvpmos >>
rect -100 483 100 683
rect -100 118 100 318
rect -100 -247 100 -47
rect -100 -612 100 -412
<< mvpdiff >>
rect -158 671 -100 683
rect -158 495 -146 671
rect -112 495 -100 671
rect -158 483 -100 495
rect 100 671 158 683
rect 100 495 112 671
rect 146 495 158 671
rect 100 483 158 495
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect -158 -59 -100 -47
rect -158 -235 -146 -59
rect -112 -235 -100 -59
rect -158 -247 -100 -235
rect 100 -59 158 -47
rect 100 -235 112 -59
rect 146 -235 158 -59
rect 100 -247 158 -235
rect -158 -424 -100 -412
rect -158 -600 -146 -424
rect -112 -600 -100 -424
rect -158 -612 -100 -600
rect 100 -424 158 -412
rect 100 -600 112 -424
rect 146 -600 158 -424
rect 100 -612 158 -600
<< mvpdiffc >>
rect -146 495 -112 671
rect 112 495 146 671
rect -146 130 -112 306
rect 112 130 146 306
rect -146 -235 -112 -59
rect 112 -235 146 -59
rect -146 -600 -112 -424
rect 112 -600 146 -424
<< mvnsubdiff >>
rect -292 831 292 843
rect -292 797 -184 831
rect 184 797 292 831
rect -292 785 292 797
rect -292 735 -234 785
rect -292 -735 -280 735
rect -246 -735 -234 735
rect 234 735 292 785
rect -292 -785 -234 -735
rect 234 -735 246 735
rect 280 -735 292 735
rect 234 -785 292 -735
rect -292 -797 292 -785
rect -292 -831 -184 -797
rect 184 -831 292 -797
rect -292 -843 292 -831
<< mvnsubdiffcont >>
rect -184 797 184 831
rect -280 -735 -246 735
rect 246 -735 280 735
rect -184 -831 184 -797
<< poly >>
rect -100 683 100 709
rect -100 436 100 483
rect -100 402 -84 436
rect 84 402 100 436
rect -100 386 100 402
rect -100 318 100 344
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -47 100 -21
rect -100 -294 100 -247
rect -100 -328 -84 -294
rect 84 -328 100 -294
rect -100 -344 100 -328
rect -100 -412 100 -386
rect -100 -659 100 -612
rect -100 -693 -84 -659
rect 84 -693 100 -659
rect -100 -709 100 -693
<< polycont >>
rect -84 402 84 436
rect -84 37 84 71
rect -84 -328 84 -294
rect -84 -693 84 -659
<< locali >>
rect -280 797 -184 831
rect 184 797 280 831
rect -280 735 -246 797
rect 246 735 280 797
rect -146 671 -112 687
rect -146 479 -112 495
rect 112 671 146 687
rect 112 479 146 495
rect -100 402 -84 436
rect 84 402 100 436
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -146 -59 -112 -43
rect -146 -251 -112 -235
rect 112 -59 146 -43
rect 112 -251 146 -235
rect -100 -328 -84 -294
rect 84 -328 100 -294
rect -146 -424 -112 -408
rect -146 -616 -112 -600
rect 112 -424 146 -408
rect 112 -616 146 -600
rect -100 -693 -84 -659
rect 84 -693 100 -659
rect -280 -797 -246 -735
rect 246 -797 280 -735
rect -280 -831 -184 -797
rect 184 -831 280 -797
<< viali >>
rect -146 495 -112 671
rect 112 495 146 671
rect -84 402 84 436
rect -146 130 -112 306
rect 112 130 146 306
rect -84 37 84 71
rect -146 -235 -112 -59
rect 112 -235 146 -59
rect -84 -328 84 -294
rect -146 -600 -112 -424
rect 112 -600 146 -424
rect -84 -693 84 -659
<< metal1 >>
rect -152 671 -106 683
rect -152 495 -146 671
rect -112 495 -106 671
rect -152 483 -106 495
rect 106 671 152 683
rect 106 495 112 671
rect 146 495 152 671
rect 106 483 152 495
rect -96 436 96 442
rect -96 402 -84 436
rect 84 402 96 436
rect -96 396 96 402
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -152 -59 -106 -47
rect -152 -235 -146 -59
rect -112 -235 -106 -59
rect -152 -247 -106 -235
rect 106 -59 152 -47
rect 106 -235 112 -59
rect 146 -235 152 -59
rect 106 -247 152 -235
rect -96 -294 96 -288
rect -96 -328 -84 -294
rect 84 -328 96 -294
rect -96 -334 96 -328
rect -152 -424 -106 -412
rect -152 -600 -146 -424
rect -112 -600 -106 -424
rect -152 -612 -106 -600
rect 106 -424 152 -412
rect 106 -600 112 -424
rect 146 -600 152 -424
rect 106 -612 152 -600
rect -96 -659 96 -653
rect -96 -693 -84 -659
rect 84 -693 96 -659
rect -96 -699 96 -693
<< properties >>
string FIXED_BBOX -263 -814 263 814
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

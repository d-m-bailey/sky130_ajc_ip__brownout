magic
tech sky130A
magscale 1 2
timestamp 1712709231
<< pwell >>
rect -1819 -12582 1819 12582
<< psubdiff >>
rect -1783 12512 -1687 12546
rect 1687 12512 1783 12546
rect -1783 12450 -1749 12512
rect 1749 12450 1783 12512
rect -1783 -12512 -1749 -12450
rect 1749 -12512 1783 -12450
rect -1783 -12546 -1687 -12512
rect 1687 -12546 1783 -12512
<< psubdiffcont >>
rect -1687 12512 1687 12546
rect -1783 -12450 -1749 12450
rect 1749 -12450 1783 12450
rect -1687 -12546 1687 -12512
<< xpolycontact >>
rect -1653 11984 -1371 12416
rect -1653 -12416 -1371 -11984
rect -1275 11984 -993 12416
rect -1275 -12416 -993 -11984
rect -897 11984 -615 12416
rect -897 -12416 -615 -11984
rect -519 11984 -237 12416
rect -519 -12416 -237 -11984
rect -141 11984 141 12416
rect -141 -12416 141 -11984
rect 237 11984 519 12416
rect 237 -12416 519 -11984
rect 615 11984 897 12416
rect 615 -12416 897 -11984
rect 993 11984 1275 12416
rect 993 -12416 1275 -11984
rect 1371 11984 1653 12416
rect 1371 -12416 1653 -11984
<< xpolyres >>
rect -1653 -11984 -1371 11984
rect -1275 -11984 -993 11984
rect -897 -11984 -615 11984
rect -519 -11984 -237 11984
rect -141 -11984 141 11984
rect 237 -11984 519 11984
rect 615 -11984 897 11984
rect 993 -11984 1275 11984
rect 1371 -11984 1653 11984
<< locali >>
rect -1783 12512 -1687 12546
rect 1687 12512 1783 12546
rect -1783 12450 -1749 12512
rect 1749 12450 1783 12512
rect -1783 -12512 -1749 -12450
rect 1749 -12512 1783 -12450
rect -1783 -12546 -1687 -12512
rect 1687 -12546 1783 -12512
<< viali >>
rect -1637 12001 -1387 12398
rect -1259 12001 -1009 12398
rect -881 12001 -631 12398
rect -503 12001 -253 12398
rect -125 12001 125 12398
rect 253 12001 503 12398
rect 631 12001 881 12398
rect 1009 12001 1259 12398
rect 1387 12001 1637 12398
rect -1637 -12398 -1387 -12001
rect -1259 -12398 -1009 -12001
rect -881 -12398 -631 -12001
rect -503 -12398 -253 -12001
rect -125 -12398 125 -12001
rect 253 -12398 503 -12001
rect 631 -12398 881 -12001
rect 1009 -12398 1259 -12001
rect 1387 -12398 1637 -12001
<< metal1 >>
rect -1643 12398 -1381 12410
rect -1643 12001 -1637 12398
rect -1387 12001 -1381 12398
rect -1643 11989 -1381 12001
rect -1265 12398 -1003 12410
rect -1265 12001 -1259 12398
rect -1009 12001 -1003 12398
rect -1265 11989 -1003 12001
rect -887 12398 -625 12410
rect -887 12001 -881 12398
rect -631 12001 -625 12398
rect -887 11989 -625 12001
rect -509 12398 -247 12410
rect -509 12001 -503 12398
rect -253 12001 -247 12398
rect -509 11989 -247 12001
rect -131 12398 131 12410
rect -131 12001 -125 12398
rect 125 12001 131 12398
rect -131 11989 131 12001
rect 247 12398 509 12410
rect 247 12001 253 12398
rect 503 12001 509 12398
rect 247 11989 509 12001
rect 625 12398 887 12410
rect 625 12001 631 12398
rect 881 12001 887 12398
rect 625 11989 887 12001
rect 1003 12398 1265 12410
rect 1003 12001 1009 12398
rect 1259 12001 1265 12398
rect 1003 11989 1265 12001
rect 1381 12398 1643 12410
rect 1381 12001 1387 12398
rect 1637 12001 1643 12398
rect 1381 11989 1643 12001
rect -1643 -12001 -1381 -11989
rect -1643 -12398 -1637 -12001
rect -1387 -12398 -1381 -12001
rect -1643 -12410 -1381 -12398
rect -1265 -12001 -1003 -11989
rect -1265 -12398 -1259 -12001
rect -1009 -12398 -1003 -12001
rect -1265 -12410 -1003 -12398
rect -887 -12001 -625 -11989
rect -887 -12398 -881 -12001
rect -631 -12398 -625 -12001
rect -887 -12410 -625 -12398
rect -509 -12001 -247 -11989
rect -509 -12398 -503 -12001
rect -253 -12398 -247 -12001
rect -509 -12410 -247 -12398
rect -131 -12001 131 -11989
rect -131 -12398 -125 -12001
rect 125 -12398 131 -12001
rect -131 -12410 131 -12398
rect 247 -12001 509 -11989
rect 247 -12398 253 -12001
rect 503 -12398 509 -12001
rect 247 -12410 509 -12398
rect 625 -12001 887 -11989
rect 625 -12398 631 -12001
rect 881 -12398 887 -12001
rect 625 -12410 887 -12398
rect 1003 -12001 1265 -11989
rect 1003 -12398 1009 -12001
rect 1259 -12398 1265 -12001
rect 1003 -12410 1265 -12398
rect 1381 -12001 1643 -11989
rect 1381 -12398 1387 -12001
rect 1637 -12398 1643 -12001
rect 1381 -12410 1643 -12398
<< properties >>
string FIXED_BBOX -1766 -12529 1766 12529
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 120 m 1 nx 9 wmin 1.410 lmin 0.50 rho 2000 val 170.479k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712901199
<< error_p >>
rect 28655 23395 28729 23469
rect 28814 22703 28888 22777
rect 29067 22024 29141 22098
<< pwell >>
rect -2026 68336 42057 68472
rect -2026 38153 -1890 68336
rect 41921 38153 42057 68336
rect -2026 38017 42057 38153
<< psubdiff >>
rect -1990 68402 -1930 68436
rect 41961 68402 42021 68436
rect -1990 68376 -1956 68402
rect -1990 38087 -1956 38113
rect 41987 68376 42021 68402
rect 41987 38087 42021 38113
rect -1990 38053 -1930 38087
rect 41961 38053 42021 38087
<< psubdiffcont >>
rect -1930 68402 41961 68436
rect -1990 38113 -1956 68376
rect 41987 38113 42021 68376
rect -1930 38053 41961 38087
<< locali >>
rect -1990 68402 -1930 68436
rect 41961 68402 42021 68436
rect -1990 68376 -1956 68402
rect -1990 38087 -1956 38113
rect 41987 68376 42021 68402
rect 41987 38087 42021 38113
rect -1990 38053 -1930 38087
rect 41961 38053 42021 38087
rect 44279 16162 44407 16290
rect 44488 16157 44552 16221
rect 44623 16162 44687 16290
rect 45359 16113 45417 16171
rect 45203 15904 45331 16032
rect 45372 15904 45436 15968
rect 45471 15904 45535 16032
rect 45317 15600 45445 15664
rect 39436 15526 39484 15574
<< viali >>
rect -1930 68402 41961 68436
rect -1990 38156 -1956 68349
rect 41987 38145 42021 68338
rect -1930 38053 41961 38087
<< metal1 >>
rect -2030 68436 42061 68476
rect -2030 68402 -1930 68436
rect 41961 68402 42061 68436
rect -2030 68349 42061 68402
rect -2030 38156 -1990 68349
rect -1956 68338 42061 68349
rect -1956 68336 41987 68338
rect -1956 38156 -1890 68336
rect -2030 38153 -1890 38156
rect 41921 38153 41987 68336
rect -2030 38145 41987 38153
rect 42021 38145 42061 68338
rect -2030 38087 42061 38145
rect -2030 38053 -1930 38087
rect 41961 38053 42061 38087
rect -2030 38013 42061 38053
<< metal3 >>
rect -2433 28873 42464 28879
rect -2433 28485 -2427 28873
rect -2039 28485 42070 28873
rect 42458 28485 42464 28873
rect -2433 28479 42464 28485
rect -2433 28413 42464 28419
rect -2433 28025 -1967 28413
rect -1579 28025 41610 28413
rect 41998 28025 42464 28413
rect -2433 28019 42464 28025
rect -2433 27953 42464 27959
rect -2433 27565 -1507 27953
rect -1119 27565 41150 27953
rect 41538 27565 42464 27953
rect -2433 27559 42464 27565
rect -2433 27493 42464 27499
rect -2433 27105 -1047 27493
rect -659 27105 40690 27493
rect 41078 27105 42464 27493
rect -2433 27099 42464 27105
rect 118 27089 528 27099
rect 28655 23395 28729 23469
rect 28814 22703 28888 22777
rect 29067 22024 29141 22098
rect -2433 -616 42464 -610
rect -2433 -1004 -1047 -616
rect -659 -1004 40690 -616
rect 41078 -1004 42464 -616
rect -2433 -1010 42464 -1004
rect -2433 -1076 42464 -1070
rect -2433 -1464 -1507 -1076
rect -1119 -1464 41150 -1076
rect 41538 -1464 42464 -1076
rect -2433 -1470 42464 -1464
rect -2433 -1536 42464 -1530
rect -2433 -1924 -1967 -1536
rect -1579 -1924 41610 -1536
rect 41998 -1924 42464 -1536
rect -2433 -1930 42464 -1924
rect -2433 -1996 42464 -1990
rect -2433 -2384 -2427 -1996
rect -2039 -2384 42070 -1996
rect 42458 -2384 42464 -1996
rect -2433 -2390 42464 -2384
<< via3 >>
rect -2427 28485 -2039 28873
rect 42070 28485 42458 28873
rect -1967 28025 -1579 28413
rect 41610 28025 41998 28413
rect -1507 27565 -1119 27953
rect 41150 27565 41538 27953
rect -1047 27105 -659 27493
rect 40690 27105 41078 27493
rect -1047 -1004 -659 -616
rect 40690 -1004 41078 -616
rect -1507 -1464 -1119 -1076
rect 41150 -1464 41538 -1076
rect -1967 -1924 -1579 -1536
rect 41610 -1924 41998 -1536
rect -2427 -2384 -2039 -1996
rect 42070 -2384 42458 -1996
<< metal4 >>
rect -2433 28873 -2033 28880
rect -2433 28485 -2427 28873
rect -2039 28485 -2033 28873
rect -2433 -1996 -2033 28485
rect -2433 -2384 -2427 -1996
rect -2039 -2384 -2033 -1996
rect -2433 -2390 -2033 -2384
rect -1973 28413 -1573 28880
rect -1973 28025 -1967 28413
rect -1579 28025 -1573 28413
rect -1973 -1536 -1573 28025
rect -1973 -1924 -1967 -1536
rect -1579 -1924 -1573 -1536
rect -1973 -2390 -1573 -1924
rect -1513 27953 -1113 28880
rect -1513 27565 -1507 27953
rect -1119 27565 -1113 27953
rect -1513 -1076 -1113 27565
rect -1513 -1464 -1507 -1076
rect -1119 -1464 -1113 -1076
rect -1513 -2390 -1113 -1464
rect -1053 27493 -653 28880
rect -1053 27105 -1047 27493
rect -659 27105 -653 27493
rect -1053 7236 -653 27105
rect 40684 27493 41084 28880
rect 40684 27105 40690 27493
rect 41078 27105 41084 27493
rect -1053 6834 -649 7236
rect -1053 -616 -653 6834
rect -1053 -1004 -1047 -616
rect -659 -1004 -653 -616
rect -1053 -2390 -653 -1004
rect 40684 -616 41084 27105
rect 40684 -1004 40690 -616
rect 41078 -1004 41084 -616
rect 40684 -2390 41084 -1004
rect 41144 27953 41544 28880
rect 41144 27565 41150 27953
rect 41538 27565 41544 27953
rect 41144 -1076 41544 27565
rect 41144 -1464 41150 -1076
rect 41538 -1464 41544 -1076
rect 41144 -2390 41544 -1464
rect 41604 28413 42004 28880
rect 41604 28025 41610 28413
rect 41998 28025 42004 28413
rect 41604 -1536 42004 28025
rect 41604 -1924 41610 -1536
rect 41998 -1924 42004 -1536
rect 41604 -2390 42004 -1924
rect 42064 28873 42464 28880
rect 42064 28485 42070 28873
rect 42458 28485 42464 28873
rect 42064 -1996 42464 28485
rect 42064 -2384 42070 -1996
rect 42458 -2384 42464 -1996
rect 42064 -2390 42464 -2384
<< labels >>
flabel metal3 894 -2390 894 -2390 0 FreeSans 1600 0 0 0 dvdd
port 3 nsew
flabel metal3 894 -1010 894 -1010 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal3 894 -1470 894 -1470 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 894 -1930 894 -1930 0 FreeSans 1600 0 0 0 dvss
port 4 nsew
<< end >>

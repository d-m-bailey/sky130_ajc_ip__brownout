magic
tech sky130A
magscale 1 2
timestamp 1712467038
<< nwell >>
rect -1653 -762 1653 762
<< mvpmos >>
rect -1395 -536 -1275 464
rect -1217 -536 -1097 464
rect -1039 -536 -919 464
rect -861 -536 -741 464
rect -683 -536 -563 464
rect -505 -536 -385 464
rect -327 -536 -207 464
rect -149 -536 -29 464
rect 29 -536 149 464
rect 207 -536 327 464
rect 385 -536 505 464
rect 563 -536 683 464
rect 741 -536 861 464
rect 919 -536 1039 464
rect 1097 -536 1217 464
rect 1275 -536 1395 464
<< mvpdiff >>
rect -1453 452 -1395 464
rect -1453 -524 -1441 452
rect -1407 -524 -1395 452
rect -1453 -536 -1395 -524
rect -1275 452 -1217 464
rect -1275 -524 -1263 452
rect -1229 -524 -1217 452
rect -1275 -536 -1217 -524
rect -1097 452 -1039 464
rect -1097 -524 -1085 452
rect -1051 -524 -1039 452
rect -1097 -536 -1039 -524
rect -919 452 -861 464
rect -919 -524 -907 452
rect -873 -524 -861 452
rect -919 -536 -861 -524
rect -741 452 -683 464
rect -741 -524 -729 452
rect -695 -524 -683 452
rect -741 -536 -683 -524
rect -563 452 -505 464
rect -563 -524 -551 452
rect -517 -524 -505 452
rect -563 -536 -505 -524
rect -385 452 -327 464
rect -385 -524 -373 452
rect -339 -524 -327 452
rect -385 -536 -327 -524
rect -207 452 -149 464
rect -207 -524 -195 452
rect -161 -524 -149 452
rect -207 -536 -149 -524
rect -29 452 29 464
rect -29 -524 -17 452
rect 17 -524 29 452
rect -29 -536 29 -524
rect 149 452 207 464
rect 149 -524 161 452
rect 195 -524 207 452
rect 149 -536 207 -524
rect 327 452 385 464
rect 327 -524 339 452
rect 373 -524 385 452
rect 327 -536 385 -524
rect 505 452 563 464
rect 505 -524 517 452
rect 551 -524 563 452
rect 505 -536 563 -524
rect 683 452 741 464
rect 683 -524 695 452
rect 729 -524 741 452
rect 683 -536 741 -524
rect 861 452 919 464
rect 861 -524 873 452
rect 907 -524 919 452
rect 861 -536 919 -524
rect 1039 452 1097 464
rect 1039 -524 1051 452
rect 1085 -524 1097 452
rect 1039 -536 1097 -524
rect 1217 452 1275 464
rect 1217 -524 1229 452
rect 1263 -524 1275 452
rect 1217 -536 1275 -524
rect 1395 452 1453 464
rect 1395 -524 1407 452
rect 1441 -524 1453 452
rect 1395 -536 1453 -524
<< mvpdiffc >>
rect -1441 -524 -1407 452
rect -1263 -524 -1229 452
rect -1085 -524 -1051 452
rect -907 -524 -873 452
rect -729 -524 -695 452
rect -551 -524 -517 452
rect -373 -524 -339 452
rect -195 -524 -161 452
rect -17 -524 17 452
rect 161 -524 195 452
rect 339 -524 373 452
rect 517 -524 551 452
rect 695 -524 729 452
rect 873 -524 907 452
rect 1051 -524 1085 452
rect 1229 -524 1263 452
rect 1407 -524 1441 452
<< mvnsubdiff >>
rect -1587 684 1587 696
rect -1587 650 -1479 684
rect 1479 650 1587 684
rect -1587 638 1587 650
rect -1587 588 -1529 638
rect -1587 -588 -1575 588
rect -1541 -588 -1529 588
rect 1529 588 1587 638
rect -1587 -638 -1529 -588
rect 1529 -588 1541 588
rect 1575 -588 1587 588
rect 1529 -638 1587 -588
rect -1587 -650 1587 -638
rect -1587 -684 -1479 -650
rect 1479 -684 1587 -650
rect -1587 -696 1587 -684
<< mvnsubdiffcont >>
rect -1479 650 1479 684
rect -1575 -588 -1541 588
rect 1541 -588 1575 588
rect -1479 -684 1479 -650
<< poly >>
rect -1395 545 -1275 561
rect -1395 511 -1379 545
rect -1291 511 -1275 545
rect -1395 464 -1275 511
rect -1217 545 -1097 561
rect -1217 511 -1201 545
rect -1113 511 -1097 545
rect -1217 464 -1097 511
rect -1039 545 -919 561
rect -1039 511 -1023 545
rect -935 511 -919 545
rect -1039 464 -919 511
rect -861 545 -741 561
rect -861 511 -845 545
rect -757 511 -741 545
rect -861 464 -741 511
rect -683 545 -563 561
rect -683 511 -667 545
rect -579 511 -563 545
rect -683 464 -563 511
rect -505 545 -385 561
rect -505 511 -489 545
rect -401 511 -385 545
rect -505 464 -385 511
rect -327 545 -207 561
rect -327 511 -311 545
rect -223 511 -207 545
rect -327 464 -207 511
rect -149 545 -29 561
rect -149 511 -133 545
rect -45 511 -29 545
rect -149 464 -29 511
rect 29 545 149 561
rect 29 511 45 545
rect 133 511 149 545
rect 29 464 149 511
rect 207 545 327 561
rect 207 511 223 545
rect 311 511 327 545
rect 207 464 327 511
rect 385 545 505 561
rect 385 511 401 545
rect 489 511 505 545
rect 385 464 505 511
rect 563 545 683 561
rect 563 511 579 545
rect 667 511 683 545
rect 563 464 683 511
rect 741 545 861 561
rect 741 511 757 545
rect 845 511 861 545
rect 741 464 861 511
rect 919 545 1039 561
rect 919 511 935 545
rect 1023 511 1039 545
rect 919 464 1039 511
rect 1097 545 1217 561
rect 1097 511 1113 545
rect 1201 511 1217 545
rect 1097 464 1217 511
rect 1275 545 1395 561
rect 1275 511 1291 545
rect 1379 511 1395 545
rect 1275 464 1395 511
rect -1395 -562 -1275 -536
rect -1217 -562 -1097 -536
rect -1039 -562 -919 -536
rect -861 -562 -741 -536
rect -683 -562 -563 -536
rect -505 -562 -385 -536
rect -327 -562 -207 -536
rect -149 -562 -29 -536
rect 29 -562 149 -536
rect 207 -562 327 -536
rect 385 -562 505 -536
rect 563 -562 683 -536
rect 741 -562 861 -536
rect 919 -562 1039 -536
rect 1097 -562 1217 -536
rect 1275 -562 1395 -536
<< polycont >>
rect -1379 511 -1291 545
rect -1201 511 -1113 545
rect -1023 511 -935 545
rect -845 511 -757 545
rect -667 511 -579 545
rect -489 511 -401 545
rect -311 511 -223 545
rect -133 511 -45 545
rect 45 511 133 545
rect 223 511 311 545
rect 401 511 489 545
rect 579 511 667 545
rect 757 511 845 545
rect 935 511 1023 545
rect 1113 511 1201 545
rect 1291 511 1379 545
<< locali >>
rect -1575 650 -1479 684
rect 1479 650 1575 684
rect -1575 588 -1541 650
rect 1541 588 1575 650
rect -1395 511 -1379 545
rect -1291 511 -1275 545
rect -1217 511 -1201 545
rect -1113 511 -1097 545
rect -1039 511 -1023 545
rect -935 511 -919 545
rect -861 511 -845 545
rect -757 511 -741 545
rect -683 511 -667 545
rect -579 511 -563 545
rect -505 511 -489 545
rect -401 511 -385 545
rect -327 511 -311 545
rect -223 511 -207 545
rect -149 511 -133 545
rect -45 511 -29 545
rect 29 511 45 545
rect 133 511 149 545
rect 207 511 223 545
rect 311 511 327 545
rect 385 511 401 545
rect 489 511 505 545
rect 563 511 579 545
rect 667 511 683 545
rect 741 511 757 545
rect 845 511 861 545
rect 919 511 935 545
rect 1023 511 1039 545
rect 1097 511 1113 545
rect 1201 511 1217 545
rect 1275 511 1291 545
rect 1379 511 1395 545
rect -1441 452 -1407 468
rect -1441 -540 -1407 -524
rect -1263 452 -1229 468
rect -1263 -540 -1229 -524
rect -1085 452 -1051 468
rect -1085 -540 -1051 -524
rect -907 452 -873 468
rect -907 -540 -873 -524
rect -729 452 -695 468
rect -729 -540 -695 -524
rect -551 452 -517 468
rect -551 -540 -517 -524
rect -373 452 -339 468
rect -373 -540 -339 -524
rect -195 452 -161 468
rect -195 -540 -161 -524
rect -17 452 17 468
rect -17 -540 17 -524
rect 161 452 195 468
rect 161 -540 195 -524
rect 339 452 373 468
rect 339 -540 373 -524
rect 517 452 551 468
rect 517 -540 551 -524
rect 695 452 729 468
rect 695 -540 729 -524
rect 873 452 907 468
rect 873 -540 907 -524
rect 1051 452 1085 468
rect 1051 -540 1085 -524
rect 1229 452 1263 468
rect 1229 -540 1263 -524
rect 1407 452 1441 468
rect 1407 -540 1441 -524
rect -1575 -650 -1541 -588
rect 1541 -650 1575 -588
rect -1575 -684 -1479 -650
rect 1479 -684 1575 -650
<< viali >>
rect -1379 511 -1291 545
rect -1201 511 -1113 545
rect -1023 511 -935 545
rect -845 511 -757 545
rect -667 511 -579 545
rect -489 511 -401 545
rect -311 511 -223 545
rect -133 511 -45 545
rect 45 511 133 545
rect 223 511 311 545
rect 401 511 489 545
rect 579 511 667 545
rect 757 511 845 545
rect 935 511 1023 545
rect 1113 511 1201 545
rect 1291 511 1379 545
rect -1441 -524 -1407 452
rect -1263 -524 -1229 452
rect -1085 -524 -1051 452
rect -907 -524 -873 452
rect -729 -524 -695 452
rect -551 -524 -517 452
rect -373 -524 -339 452
rect -195 -524 -161 452
rect -17 -524 17 452
rect 161 -524 195 452
rect 339 -524 373 452
rect 517 -524 551 452
rect 695 -524 729 452
rect 873 -524 907 452
rect 1051 -524 1085 452
rect 1229 -524 1263 452
rect 1407 -524 1441 452
<< metal1 >>
rect -1391 545 -1279 551
rect -1391 511 -1379 545
rect -1291 511 -1279 545
rect -1391 505 -1279 511
rect -1213 545 -1101 551
rect -1213 511 -1201 545
rect -1113 511 -1101 545
rect -1213 505 -1101 511
rect -1035 545 -923 551
rect -1035 511 -1023 545
rect -935 511 -923 545
rect -1035 505 -923 511
rect -857 545 -745 551
rect -857 511 -845 545
rect -757 511 -745 545
rect -857 505 -745 511
rect -679 545 -567 551
rect -679 511 -667 545
rect -579 511 -567 545
rect -679 505 -567 511
rect -501 545 -389 551
rect -501 511 -489 545
rect -401 511 -389 545
rect -501 505 -389 511
rect -323 545 -211 551
rect -323 511 -311 545
rect -223 511 -211 545
rect -323 505 -211 511
rect -145 545 -33 551
rect -145 511 -133 545
rect -45 511 -33 545
rect -145 505 -33 511
rect 33 545 145 551
rect 33 511 45 545
rect 133 511 145 545
rect 33 505 145 511
rect 211 545 323 551
rect 211 511 223 545
rect 311 511 323 545
rect 211 505 323 511
rect 389 545 501 551
rect 389 511 401 545
rect 489 511 501 545
rect 389 505 501 511
rect 567 545 679 551
rect 567 511 579 545
rect 667 511 679 545
rect 567 505 679 511
rect 745 545 857 551
rect 745 511 757 545
rect 845 511 857 545
rect 745 505 857 511
rect 923 545 1035 551
rect 923 511 935 545
rect 1023 511 1035 545
rect 923 505 1035 511
rect 1101 545 1213 551
rect 1101 511 1113 545
rect 1201 511 1213 545
rect 1101 505 1213 511
rect 1279 545 1391 551
rect 1279 511 1291 545
rect 1379 511 1391 545
rect 1279 505 1391 511
rect -1447 452 -1401 464
rect -1447 -524 -1441 452
rect -1407 -524 -1401 452
rect -1447 -536 -1401 -524
rect -1269 452 -1223 464
rect -1269 -524 -1263 452
rect -1229 -524 -1223 452
rect -1269 -536 -1223 -524
rect -1091 452 -1045 464
rect -1091 -524 -1085 452
rect -1051 -524 -1045 452
rect -1091 -536 -1045 -524
rect -913 452 -867 464
rect -913 -524 -907 452
rect -873 -524 -867 452
rect -913 -536 -867 -524
rect -735 452 -689 464
rect -735 -524 -729 452
rect -695 -524 -689 452
rect -735 -536 -689 -524
rect -557 452 -511 464
rect -557 -524 -551 452
rect -517 -524 -511 452
rect -557 -536 -511 -524
rect -379 452 -333 464
rect -379 -524 -373 452
rect -339 -524 -333 452
rect -379 -536 -333 -524
rect -201 452 -155 464
rect -201 -524 -195 452
rect -161 -524 -155 452
rect -201 -536 -155 -524
rect -23 452 23 464
rect -23 -524 -17 452
rect 17 -524 23 452
rect -23 -536 23 -524
rect 155 452 201 464
rect 155 -524 161 452
rect 195 -524 201 452
rect 155 -536 201 -524
rect 333 452 379 464
rect 333 -524 339 452
rect 373 -524 379 452
rect 333 -536 379 -524
rect 511 452 557 464
rect 511 -524 517 452
rect 551 -524 557 452
rect 511 -536 557 -524
rect 689 452 735 464
rect 689 -524 695 452
rect 729 -524 735 452
rect 689 -536 735 -524
rect 867 452 913 464
rect 867 -524 873 452
rect 907 -524 913 452
rect 867 -536 913 -524
rect 1045 452 1091 464
rect 1045 -524 1051 452
rect 1085 -524 1091 452
rect 1045 -536 1091 -524
rect 1223 452 1269 464
rect 1223 -524 1229 452
rect 1263 -524 1269 452
rect 1223 -536 1269 -524
rect 1401 452 1447 464
rect 1401 -524 1407 452
rect 1441 -524 1447 452
rect 1401 -536 1447 -524
<< properties >>
string FIXED_BBOX -1558 -667 1558 667
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

* NGSPICE file created from brownout_dig.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

.subckt brownout_dig VGND VPWR brout_filt ena force_rc_osc force_short_oneshot osc_ck
+ osc_ck_256 osc_ena otrip[0] otrip[1] otrip[2] otrip_decoded[0] otrip_decoded[1]
+ otrip_decoded[2] otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6]
+ otrip_decoded[7] out_unbuf timed_out vtrip[0] vtrip[1] vtrip[2] vtrip_decoded[0]
+ vtrip_decoded[1] vtrip_decoded[2] vtrip_decoded[3] vtrip_decoded[4] vtrip_decoded[5]
+ vtrip_decoded[6] vtrip_decoded[7]
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_131_ net10 net9 net8 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__and3b_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_114_ _063_ _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput20 net20 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ net10 net8 net9 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__nor3b_1
XFILLER_0_19_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_113_ cnt\[5\] cnt\[6\] VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__and2_1
Xclkbuf_2_3__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_3__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR out_unbuf sky130_fd_sc_hd__buf_2
XFILLER_0_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_112_ cnt\[4\] _062_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__and2_1
Xhold10 _001_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput11 net11 VGND VGND VPWR VPWR osc_ck_256 sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR timed_out sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ clknet_2_1__leaf_osc_ck net41 brout_filt_ena_rsb VGND VGND VPWR VPWR brout_filt_retime_rsb
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_111_ cnt\[1\] cnt\[0\] cnt\[3\] cnt\[2\] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold11 cnt_ck_256\[0\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR vtrip_decoded[0] sky130_fd_sc_hd__buf_2
XFILLER_0_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_187_ clknet_2_1__leaf_osc_ck net37 brout_filt_ena_rsb VGND VGND VPWR VPWR brout_filt_retime_rsb_stg1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nand2_1
Xhold12 cnt_ck_256\[2\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__clkbuf_4
Xoutput24 net24 VGND VGND VPWR VPWR vtrip_decoded[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_186_ clknet_2_1__leaf_osc_ck net39 net38 VGND VGND VPWR VPWR brout_filt_retimed
+ sky130_fd_sc_hd__dfrtp_1
X_169_ clknet_2_2__leaf_osc_ck _018_ net35 VGND VGND VPWR VPWR cnt\[11\] sky130_fd_sc_hd__dfstp_1
Xhold13 cnt_ck_256\[4\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_11_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR vtrip_decoded[2] sky130_fd_sc_hd__buf_2
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_185_ clknet_2_1__leaf_osc_ck net1 net38 VGND VGND VPWR VPWR brout_filt_retimed_stg1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_168_ clknet_2_2__leaf_osc_ck _017_ net34 VGND VGND VPWR VPWR cnt\[10\] sky130_fd_sc_hd__dfstp_1
X_099_ cnt\[12\] _053_ net53 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a21oi_1
Xhold14 cnt_ck_256\[5\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR vtrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ clknet_2_0__leaf_osc_ck net42 net2 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
X_167_ clknet_2_2__leaf_osc_ck _016_ net34 VGND VGND VPWR VPWR cnt\[9\] sky130_fd_sc_hd__dfstp_1
X_098_ net33 _054_ _025_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 cnt_ck_256\[3\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR vtrip_decoded[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_182__36 VGND VGND VPWR VPWR net36 _182__36/LO sky130_fd_sc_hd__conb_1
XFILLER_0_4_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_183_ clknet_2_0__leaf_osc_ck net40 net2 VGND VGND VPWR VPWR cnt_rsb_stg2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_166_ clknet_2_2__leaf_osc_ck _015_ net34 VGND VGND VPWR VPWR cnt\[8\] sky130_fd_sc_hd__dfstp_1
X_097_ cnt\[12\] _053_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 cnt\[13\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
X_149_ net50 _028_ net51 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a21oi_1
Xoutput28 net28 VGND VGND VPWR VPWR vtrip_decoded[5] sky130_fd_sc_hd__buf_2
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ clknet_2_0__leaf_osc_ck net36 net2 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_096_ _066_ _067_ net4 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a21o_1
X_165_ clknet_2_0__leaf_osc_ck _014_ net34 VGND VGND VPWR VPWR cnt\[7\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_19_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold17 cnt\[15\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
X_148_ cnt_ck_256\[5\] cnt_ck_256\[4\] _028_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
X_079_ net31 _042_ net32 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a21oi_1
Xoutput29 net29 VGND VGND VPWR VPWR vtrip_decoded[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_2__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_181_ clknet_2_3__leaf_osc_ck net45 net38 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout31 _034_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_095_ net31 _052_ net33 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21oi_1
X_164_ clknet_2_0__leaf_osc_ck _013_ net34 VGND VGND VPWR VPWR cnt\[6\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_10_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold18 cnt_ck_256\[6\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
X_078_ cnt\[5\] _063_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_147_ net50 _028_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__xor2_1
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout32 brout_filt_retimed VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
X_180_ clknet_2_3__leaf_osc_ck _006_ net38 VGND VGND VPWR VPWR cnt_ck_256\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_094_ cnt\[11\] _049_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__xnor2_1
X_163_ clknet_2_0__leaf_osc_ck _012_ net34 VGND VGND VPWR VPWR cnt\[5\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_10_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_146_ _028_ _029_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nor2_1
X_077_ net31 _041_ net32 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_129_ net10 net9 net8 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nor3b_1
Xfanout33 brout_filt_retimed VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
X_093_ net31 _051_ net33 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a21oi_1
X_162_ clknet_2_0__leaf_osc_ck _011_ net34 VGND VGND VPWR VPWR cnt\[4\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_7_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 brout_filt VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ _063_ _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__or2_1
X_145_ net52 _026_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_128_ net10 net9 net8 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__nor3_1
XFILLER_0_17_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout34 net43 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_161_ clknet_2_0__leaf_osc_ck _010_ net34 VGND VGND VPWR VPWR cnt\[3\] sky130_fd_sc_hd__dfstp_1
X_092_ _049_ _050_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nand2b_1
Xinput2 ena VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_144_ cnt_ck_256\[3\] _026_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ cnt\[4\] _062_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nor2_1
X_127_ net7 net5 net6 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_10_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout35 net43 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_091_ cnt\[9\] cnt\[8\] _066_ cnt\[10\] VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a31o_1
X_160_ clknet_2_3__leaf_osc_ck _009_ net35 VGND VGND VPWR VPWR cnt\[2\] sky130_fd_sc_hd__dfstp_1
Xinput3 force_rc_osc VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_143_ _026_ _027_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor2_1
X_074_ net31 _039_ net32 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_126_ net5 net6 net7 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and3b_1
XFILLER_0_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ net48 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ cnt\[9\] cnt\[8\] cnt\[10\] _066_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__and4_1
Xinput4 force_short_oneshot VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ cnt_ck_256\[0\] net46 net49 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_073_ _062_ _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_125_ net6 net5 net7 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and3b_1
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_108_ net44 _032_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 otrip[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_141_ cnt_ck_256\[0\] cnt_ck_256\[1\] cnt_ck_256\[2\] VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and3_1
X_072_ cnt\[1\] cnt\[0\] cnt\[2\] cnt\[3\] VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_124_ net5 net6 net7 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__nor3b_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ net33 _059_ _060_ _025_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_14_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 otrip[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_2_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_071_ _034_ _037_ net32 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_140_ cnt_ck_256\[0\] net46 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ net7 net5 net6 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and3b_1
XFILLER_0_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_106_ cnt\[15\] _068_ _053_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 otrip[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_070_ cnt\[2\] _061_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_122_ net7 net5 net6 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 vtrip[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_2_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_105_ _068_ _053_ net54 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 vtrip[0] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ net7 net6 net5 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__nor3b_1
X_104_ _057_ _058_ net21 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 vtrip[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ net7 net5 net6 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_6_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_103_ _068_ _053_ net33 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 brout_filt_retime_rsb VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_179_ clknet_2_3__leaf_osc_ck _005_ net38 VGND VGND VPWR VPWR cnt_ck_256\[5\] sky130_fd_sc_hd__dfrtp_1
X_102_ cnt\[13\] cnt\[12\] _053_ cnt\[14\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__a31o_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 brout_filt_retimed_stg1 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_178_ clknet_2_3__leaf_osc_ck _004_ net38 VGND VGND VPWR VPWR cnt_ck_256\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_101_ _055_ _056_ _025_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 cnt_rsb_stg1 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_177_ clknet_2_1__leaf_osc_ck _003_ net38 VGND VGND VPWR VPWR cnt_ck_256\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_100_ cnt\[13\] cnt\[12\] _053_ net33 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 brout_filt_retime_rsb_stg1 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_176_ clknet_2_1__leaf_osc_ck _002_ net38 VGND VGND VPWR VPWR cnt_ck_256\[2\] sky130_fd_sc_hd__dfrtp_1
X_159_ clknet_2_3__leaf_osc_ck _008_ net35 VGND VGND VPWR VPWR cnt\[1\] sky130_fd_sc_hd__dfstp_1
Xhold5 cnt_rsb_stg2 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_187__37 VGND VGND VPWR VPWR net37 _187__37/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_11_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_175_ clknet_2_1__leaf_osc_ck net47 net38 VGND VGND VPWR VPWR cnt_ck_256\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ net31 _048_ net32 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a21oi_1
X_158_ clknet_2_0__leaf_osc_ck _007_ net34 VGND VGND VPWR VPWR cnt\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 cnt_rsb VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_174_ clknet_2_1__leaf_osc_ck _000_ net38 VGND VGND VPWR VPWR cnt_ck_256\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_088_ cnt\[9\] _046_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__xor2_1
X_157_ _061_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 net11 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_7_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_173_ clknet_2_2__leaf_osc_ck _022_ net35 VGND VGND VPWR VPWR cnt\[15\] sky130_fd_sc_hd__dfstp_1
X_087_ net31 _047_ net32 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a21oi_1
X_156_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 _023_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
X_139_ net2 _025_ brout_filt_ena_rsb net3 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_17_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_172_ clknet_2_2__leaf_osc_ck _021_ net35 VGND VGND VPWR VPWR cnt\[14\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_5_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_086_ cnt\[8\] _066_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__xnor2_1
X_155_ cnt\[0\] net31 net32 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21oi_1
Xhold9 cnt_ck_256\[1\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
X_069_ _034_ _036_ net32 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21oi_1
X_138_ net1 net2 VGND VGND VPWR VPWR brout_filt_ena_rsb sky130_fd_sc_hd__and2_1
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_171_ clknet_2_2__leaf_osc_ck _020_ net35 VGND VGND VPWR VPWR cnt\[13\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_154_ net4 net22 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ cnt\[8\] _066_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_137_ net33 _024_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ clknet_2_2__leaf_osc_ck _019_ net34 VGND VGND VPWR VPWR cnt\[12\] sky130_fd_sc_hd__dfstp_1
X_084_ net31 _045_ net32 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ _032_ _033_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and2_1
X_136_ cnt\[15\] _066_ _067_ _068_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_119_ net33 net22 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and2b_1
XFILLER_0_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ cnt\[7\] _065_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__xor2_1
X_152_ net55 _030_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ net10 net9 net8 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__and3_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_118_ cnt\[15\] _066_ _067_ _068_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__and4_1
XFILLER_0_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_151_ cnt_ck_256\[6\] _030_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand2_1
X_082_ net31 _044_ net32 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_134_ net8 net9 net10 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__and3b_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ cnt\[13\] cnt\[12\] cnt\[14\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_12_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_081_ _065_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_0_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_150_ _030_ _031_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_133_ net9 net8 net10 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__and3b_1
XFILLER_0_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_116_ cnt\[9\] cnt\[8\] cnt\[11\] cnt\[10\] VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_20_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_080_ cnt\[5\] cnt\[4\] _062_ cnt\[6\] VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_132_ net9 net8 net10 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__nor3b_1
XFILLER_0_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_115_ cnt\[4\] cnt\[7\] _062_ _064_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_20_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput30 net30 VGND VGND VPWR VPWR vtrip_decoded[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends


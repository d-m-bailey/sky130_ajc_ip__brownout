magic
tech sky130A
magscale 1 2
timestamp 1712846855
<< pwell >>
rect -2008 -11082 2008 11082
<< psubdiff >>
rect -1972 11012 -1876 11046
rect 1876 11012 1972 11046
rect -1972 10950 -1938 11012
rect 1938 10950 1972 11012
rect -1972 -11012 -1938 -10950
rect 1938 -11012 1972 -10950
rect -1972 -11046 -1876 -11012
rect 1876 -11046 1972 -11012
<< psubdiffcont >>
rect -1876 11012 1876 11046
rect -1972 -10950 -1938 10950
rect 1938 -10950 1972 10950
rect -1876 -11046 1876 -11012
<< xpolycontact >>
rect -1842 10484 -1560 10916
rect -1842 -10916 -1560 -10484
rect -1464 10484 -1182 10916
rect -1464 -10916 -1182 -10484
rect -1086 10484 -804 10916
rect -1086 -10916 -804 -10484
rect -708 10484 -426 10916
rect -708 -10916 -426 -10484
rect -330 10484 -48 10916
rect -330 -10916 -48 -10484
rect 48 10484 330 10916
rect 48 -10916 330 -10484
rect 426 10484 708 10916
rect 426 -10916 708 -10484
rect 804 10484 1086 10916
rect 804 -10916 1086 -10484
rect 1182 10484 1464 10916
rect 1182 -10916 1464 -10484
rect 1560 10484 1842 10916
rect 1560 -10916 1842 -10484
<< xpolyres >>
rect -1842 -10484 -1560 10484
rect -1464 -10484 -1182 10484
rect -1086 -10484 -804 10484
rect -708 -10484 -426 10484
rect -330 -10484 -48 10484
rect 48 -10484 330 10484
rect 426 -10484 708 10484
rect 804 -10484 1086 10484
rect 1182 -10484 1464 10484
rect 1560 -10484 1842 10484
<< locali >>
rect -1972 11012 -1876 11046
rect 1876 11012 1972 11046
rect -1972 10950 -1938 11012
rect 1938 10950 1972 11012
rect -1972 -11012 -1938 -10950
rect 1938 -11012 1972 -10950
rect -1972 -11046 -1876 -11012
rect 1876 -11046 1972 -11012
<< viali >>
rect -1826 10501 -1576 10898
rect -1448 10501 -1198 10898
rect -1070 10501 -820 10898
rect -692 10501 -442 10898
rect -314 10501 -64 10898
rect 64 10501 314 10898
rect 442 10501 692 10898
rect 820 10501 1070 10898
rect 1198 10501 1448 10898
rect 1576 10501 1826 10898
rect -1826 -10898 -1576 -10501
rect -1448 -10898 -1198 -10501
rect -1070 -10898 -820 -10501
rect -692 -10898 -442 -10501
rect -314 -10898 -64 -10501
rect 64 -10898 314 -10501
rect 442 -10898 692 -10501
rect 820 -10898 1070 -10501
rect 1198 -10898 1448 -10501
rect 1576 -10898 1826 -10501
<< metal1 >>
rect -1832 10898 -1570 10910
rect -1832 10501 -1826 10898
rect -1576 10501 -1570 10898
rect -1832 10489 -1570 10501
rect -1454 10898 -1192 10910
rect -1454 10501 -1448 10898
rect -1198 10501 -1192 10898
rect -1454 10489 -1192 10501
rect -1076 10898 -814 10910
rect -1076 10501 -1070 10898
rect -820 10501 -814 10898
rect -1076 10489 -814 10501
rect -698 10898 -436 10910
rect -698 10501 -692 10898
rect -442 10501 -436 10898
rect -698 10489 -436 10501
rect -320 10898 -58 10910
rect -320 10501 -314 10898
rect -64 10501 -58 10898
rect -320 10489 -58 10501
rect 58 10898 320 10910
rect 58 10501 64 10898
rect 314 10501 320 10898
rect 58 10489 320 10501
rect 436 10898 698 10910
rect 436 10501 442 10898
rect 692 10501 698 10898
rect 436 10489 698 10501
rect 814 10898 1076 10910
rect 814 10501 820 10898
rect 1070 10501 1076 10898
rect 814 10489 1076 10501
rect 1192 10898 1454 10910
rect 1192 10501 1198 10898
rect 1448 10501 1454 10898
rect 1192 10489 1454 10501
rect 1570 10898 1832 10910
rect 1570 10501 1576 10898
rect 1826 10501 1832 10898
rect 1570 10489 1832 10501
rect -1832 -10501 -1570 -10489
rect -1832 -10898 -1826 -10501
rect -1576 -10898 -1570 -10501
rect -1832 -10910 -1570 -10898
rect -1454 -10501 -1192 -10489
rect -1454 -10898 -1448 -10501
rect -1198 -10898 -1192 -10501
rect -1454 -10910 -1192 -10898
rect -1076 -10501 -814 -10489
rect -1076 -10898 -1070 -10501
rect -820 -10898 -814 -10501
rect -1076 -10910 -814 -10898
rect -698 -10501 -436 -10489
rect -698 -10898 -692 -10501
rect -442 -10898 -436 -10501
rect -698 -10910 -436 -10898
rect -320 -10501 -58 -10489
rect -320 -10898 -314 -10501
rect -64 -10898 -58 -10501
rect -320 -10910 -58 -10898
rect 58 -10501 320 -10489
rect 58 -10898 64 -10501
rect 314 -10898 320 -10501
rect 58 -10910 320 -10898
rect 436 -10501 698 -10489
rect 436 -10898 442 -10501
rect 692 -10898 698 -10501
rect 436 -10910 698 -10898
rect 814 -10501 1076 -10489
rect 814 -10898 820 -10501
rect 1070 -10898 1076 -10501
rect 814 -10910 1076 -10898
rect 1192 -10501 1454 -10489
rect 1192 -10898 1198 -10501
rect 1448 -10898 1454 -10501
rect 1192 -10910 1454 -10898
rect 1570 -10501 1832 -10489
rect 1570 -10898 1576 -10501
rect 1826 -10898 1832 -10501
rect 1570 -10910 1832 -10898
<< properties >>
string FIXED_BBOX -1955 -11029 1955 11029
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 105 m 1 nx 10 wmin 1.410 lmin 0.50 rho 2000 val 149.203k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713147927
<< viali >>
rect 4169 10761 4203 10795
rect 4813 10761 4847 10795
rect 5365 10761 5399 10795
rect 5917 10761 5951 10795
rect 6745 10761 6779 10795
rect 7297 10761 7331 10795
rect 1777 10625 1811 10659
rect 2697 10625 2731 10659
rect 4077 10625 4111 10659
rect 4721 10625 4755 10659
rect 5273 10625 5307 10659
rect 5825 10625 5859 10659
rect 6653 10625 6687 10659
rect 7573 10625 7607 10659
rect 7941 10625 7975 10659
rect 2053 10557 2087 10591
rect 2973 10557 3007 10591
rect 8217 10557 8251 10591
rect 2697 10217 2731 10251
rect 3617 10217 3651 10251
rect 4997 10217 5031 10251
rect 5457 10217 5491 10251
rect 5641 10217 5675 10251
rect 6101 10217 6135 10251
rect 6285 10217 6319 10251
rect 6745 10217 6779 10251
rect 7205 10217 7239 10251
rect 7389 10217 7423 10251
rect 8033 10217 8067 10251
rect 4905 10149 4939 10183
rect 5733 10149 5767 10183
rect 6929 10149 6963 10183
rect 3341 10081 3375 10115
rect 4261 10081 4295 10115
rect 4353 10081 4387 10115
rect 4445 10081 4479 10115
rect 4629 10081 4663 10115
rect 3249 10013 3283 10047
rect 3433 10013 3467 10047
rect 4997 10013 5031 10047
rect 5089 10013 5123 10047
rect 6377 10013 6411 10047
rect 2973 9945 3007 9979
rect 4721 9945 4755 9979
rect 7021 9945 7055 9979
rect 7941 9945 7975 9979
rect 5457 9877 5491 9911
rect 6101 9877 6135 9911
rect 6745 9877 6779 9911
rect 7231 9877 7265 9911
rect 3433 9673 3467 9707
rect 3709 9537 3743 9571
rect 3801 9537 3835 9571
rect 3617 9469 3651 9503
rect 4721 9129 4755 9163
rect 3249 9061 3283 9095
rect 1685 8925 1719 8959
rect 3525 8925 3559 8959
rect 6285 8925 6319 8959
rect 6653 8925 6687 8959
rect 6929 8925 6963 8959
rect 7297 8925 7331 8959
rect 1501 8857 1535 8891
rect 3249 8857 3283 8891
rect 4169 8857 4203 8891
rect 4353 8857 4387 8891
rect 4537 8857 4571 8891
rect 3433 8789 3467 8823
rect 4077 8789 4111 8823
rect 4859 8789 4893 8823
rect 8723 8789 8757 8823
rect 5174 8585 5208 8619
rect 8861 8585 8895 8619
rect 6653 8517 6687 8551
rect 7205 8517 7239 8551
rect 2697 8449 2731 8483
rect 4537 8449 4571 8483
rect 4997 8449 5031 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5818 8449 5852 8483
rect 6469 8449 6503 8483
rect 6745 8449 6779 8483
rect 7849 8449 7883 8483
rect 7941 8449 7975 8483
rect 8401 8449 8435 8483
rect 9045 8449 9079 8483
rect 9321 8449 9355 8483
rect 9413 8449 9447 8483
rect 2329 8381 2363 8415
rect 4629 8381 4663 8415
rect 4905 8381 4939 8415
rect 7481 8381 7515 8415
rect 8493 8381 8527 8415
rect 5457 8313 5491 8347
rect 6837 8313 6871 8347
rect 8769 8313 8803 8347
rect 9229 8313 9263 8347
rect 9597 8313 9631 8347
rect 4123 8245 4157 8279
rect 5733 8245 5767 8279
rect 6469 8245 6503 8279
rect 7205 8245 7239 8279
rect 7389 8245 7423 8279
rect 7665 8245 7699 8279
rect 5411 8041 5445 8075
rect 8677 8041 8711 8075
rect 5273 7973 5307 8007
rect 7573 7973 7607 8007
rect 7665 7973 7699 8007
rect 9505 7973 9539 8007
rect 1777 7905 1811 7939
rect 4445 7905 4479 7939
rect 7205 7905 7239 7939
rect 8953 7905 8987 7939
rect 2145 7837 2179 7871
rect 3571 7837 3605 7871
rect 4997 7837 5031 7871
rect 6837 7837 6871 7871
rect 7297 7837 7331 7871
rect 7481 7837 7515 7871
rect 7757 7837 7791 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 8355 7837 8389 7871
rect 8585 7837 8619 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9689 7837 9723 7871
rect 4721 7769 4755 7803
rect 8217 7769 8251 7803
rect 3801 7701 3835 7735
rect 4905 7701 4939 7735
rect 5089 7701 5123 7735
rect 8493 7701 8527 7735
rect 9321 7701 9355 7735
rect 3157 7497 3191 7531
rect 6469 7497 6503 7531
rect 6837 7497 6871 7531
rect 7113 7497 7147 7531
rect 7297 7497 7331 7531
rect 9643 7497 9677 7531
rect 3525 7429 3559 7463
rect 7481 7429 7515 7463
rect 2973 7361 3007 7395
rect 3249 7361 3283 7395
rect 3341 7361 3375 7395
rect 3617 7361 3651 7395
rect 3709 7361 3743 7395
rect 6377 7361 6411 7395
rect 6653 7361 6687 7395
rect 7205 7361 7239 7395
rect 8217 7361 8251 7395
rect 4077 7293 4111 7327
rect 7849 7293 7883 7327
rect 2973 7225 3007 7259
rect 3341 7225 3375 7259
rect 6929 7225 6963 7259
rect 5503 7157 5537 7191
rect 8309 6953 8343 6987
rect 8953 6953 8987 6987
rect 4169 6817 4203 6851
rect 4353 6817 4387 6851
rect 4445 6817 4479 6851
rect 9321 6817 9355 6851
rect 3525 6749 3559 6783
rect 3617 6749 3651 6783
rect 4261 6749 4295 6783
rect 5089 6749 5123 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 3341 6681 3375 6715
rect 7021 6681 7055 6715
rect 3439 6613 3473 6647
rect 4629 6613 4663 6647
rect 6377 6613 6411 6647
rect 9597 6613 9631 6647
rect 4997 6409 5031 6443
rect 5641 6409 5675 6443
rect 9413 6409 9447 6443
rect 4859 6341 4893 6375
rect 3065 6273 3099 6307
rect 3433 6273 3467 6307
rect 5211 6273 5245 6307
rect 5365 6273 5399 6307
rect 5457 6273 5491 6307
rect 5825 6273 5859 6307
rect 6009 6273 6043 6307
rect 6561 6273 6595 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 8677 6273 8711 6307
rect 9689 6273 9723 6307
rect 6469 6205 6503 6239
rect 8493 6205 8527 6239
rect 8953 6205 8987 6239
rect 6929 6137 6963 6171
rect 7297 6137 7331 6171
rect 9229 6137 9263 6171
rect 2237 6069 2271 6103
rect 5825 6069 5859 6103
rect 8861 6069 8895 6103
rect 9505 6069 9539 6103
rect 3893 5865 3927 5899
rect 4353 5865 4387 5899
rect 5365 5865 5399 5899
rect 6699 5865 6733 5899
rect 9045 5865 9079 5899
rect 4813 5797 4847 5831
rect 1777 5729 1811 5763
rect 6101 5729 6135 5763
rect 8493 5729 8527 5763
rect 9229 5729 9263 5763
rect 2145 5661 2179 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 5457 5661 5491 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 8125 5661 8159 5695
rect 8585 5661 8619 5695
rect 8953 5661 8987 5695
rect 5089 5593 5123 5627
rect 5181 5593 5215 5627
rect 1593 5525 1627 5559
rect 3571 5525 3605 5559
rect 4997 5525 5031 5559
rect 6469 5525 6503 5559
rect 8769 5525 8803 5559
rect 9505 5525 9539 5559
rect 2789 5321 2823 5355
rect 3157 5321 3191 5355
rect 4997 5321 5031 5355
rect 7113 5321 7147 5355
rect 7481 5321 7515 5355
rect 9689 5321 9723 5355
rect 4629 5253 4663 5287
rect 7297 5253 7331 5287
rect 7665 5253 7699 5287
rect 8217 5253 8251 5287
rect 4813 5185 4847 5219
rect 5089 5185 5123 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 5549 5185 5583 5219
rect 5641 5185 5675 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 6561 5185 6595 5219
rect 7021 5185 7055 5219
rect 7389 5185 7423 5219
rect 2145 5117 2179 5151
rect 5825 5117 5859 5151
rect 6469 5117 6503 5151
rect 6929 5117 6963 5151
rect 7941 5117 7975 5151
rect 7297 5049 7331 5083
rect 4813 4981 4847 5015
rect 5181 4981 5215 5015
rect 7665 4981 7699 5015
rect 1409 4777 1443 4811
rect 6515 4777 6549 4811
rect 3341 4709 3375 4743
rect 6791 4709 6825 4743
rect 3157 4641 3191 4675
rect 4721 4641 4755 4675
rect 5089 4641 5123 4675
rect 8585 4641 8619 4675
rect 9045 4641 9079 4675
rect 9321 4641 9355 4675
rect 3341 4573 3375 4607
rect 3525 4573 3559 4607
rect 3617 4573 3651 4607
rect 4445 4573 4479 4607
rect 8217 4573 8251 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 2881 4505 2915 4539
rect 3801 4505 3835 4539
rect 9505 4437 9539 4471
rect 2145 4233 2179 4267
rect 5365 4233 5399 4267
rect 9229 4233 9263 4267
rect 1409 4097 1443 4131
rect 2237 4097 2271 4131
rect 2329 4097 2363 4131
rect 3157 4097 3191 4131
rect 3525 4097 3559 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 8861 4097 8895 4131
rect 9137 4097 9171 4131
rect 9413 4097 9447 4131
rect 4951 4029 4985 4063
rect 1593 3961 1627 3995
rect 9045 3961 9079 3995
rect 2421 3893 2455 3927
rect 9597 3893 9631 3927
rect 4077 3689 4111 3723
rect 3157 3621 3191 3655
rect 1409 3553 1443 3587
rect 4445 3553 4479 3587
rect 4353 3485 4387 3519
rect 7757 3485 7791 3519
rect 7849 3485 7883 3519
rect 1685 3417 1719 3451
rect 7573 3417 7607 3451
rect 7849 3349 7883 3383
rect 7573 3145 7607 3179
rect 6929 3077 6963 3111
rect 8217 3077 8251 3111
rect 8645 3077 8679 3111
rect 8861 3077 8895 3111
rect 4445 3009 4479 3043
rect 4813 3009 4847 3043
rect 4997 3009 5031 3043
rect 6009 3009 6043 3043
rect 6561 3009 6595 3043
rect 7849 3009 7883 3043
rect 9413 3009 9447 3043
rect 4261 2941 4295 2975
rect 4353 2941 4387 2975
rect 4905 2941 4939 2975
rect 5825 2941 5859 2975
rect 5917 2941 5951 2975
rect 6193 2941 6227 2975
rect 7205 2873 7239 2907
rect 4077 2805 4111 2839
rect 4629 2805 4663 2839
rect 6929 2805 6963 2839
rect 7113 2805 7147 2839
rect 7573 2805 7607 2839
rect 7757 2805 7791 2839
rect 8217 2805 8251 2839
rect 8401 2805 8435 2839
rect 8493 2805 8527 2839
rect 8677 2805 8711 2839
rect 9597 2805 9631 2839
rect 7849 2533 7883 2567
rect 4077 2465 4111 2499
rect 5549 2465 5583 2499
rect 6653 2465 6687 2499
rect 3617 2397 3651 2431
rect 3801 2397 3835 2431
rect 4721 2397 4755 2431
rect 5273 2397 5307 2431
rect 6377 2397 6411 2431
rect 7297 2397 7331 2431
rect 7665 2397 7699 2431
rect 8033 2397 8067 2431
rect 8493 2397 8527 2431
rect 9137 2397 9171 2431
rect 3433 2261 3467 2295
rect 4905 2261 4939 2295
rect 7481 2261 7515 2295
rect 8217 2261 8251 2295
rect 8677 2261 8711 2295
rect 9321 2261 9355 2295
<< metal1 >>
rect 1104 10906 10028 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 10028 10906
rect 1104 10832 10028 10854
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 3936 10764 4169 10792
rect 3936 10752 3942 10764
rect 4157 10761 4169 10764
rect 4203 10761 4215 10795
rect 4157 10755 4215 10761
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4580 10764 4813 10792
rect 4580 10752 4586 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5353 10795 5411 10801
rect 5353 10792 5365 10795
rect 5316 10764 5365 10792
rect 5316 10752 5322 10764
rect 5353 10761 5365 10764
rect 5399 10761 5411 10795
rect 5353 10755 5411 10761
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 5905 10795 5963 10801
rect 5905 10792 5917 10795
rect 5868 10764 5917 10792
rect 5868 10752 5874 10764
rect 5905 10761 5917 10764
rect 5951 10761 5963 10795
rect 5905 10755 5963 10761
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 6512 10764 6745 10792
rect 6512 10752 6518 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7156 10764 7297 10792
rect 7156 10752 7162 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1946 10656 1952 10668
rect 1811 10628 1952 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2648 10628 2697 10656
rect 2648 10616 2654 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 4062 10616 4068 10668
rect 4120 10616 4126 10668
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4672 10628 4721 10656
rect 4672 10616 4678 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 5258 10616 5264 10668
rect 5316 10616 5322 10668
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8386 10656 8392 10668
rect 7975 10628 8392 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 2038 10548 2044 10600
rect 2096 10548 2102 10600
rect 2958 10548 2964 10600
rect 3016 10548 3022 10600
rect 8202 10548 8208 10600
rect 8260 10548 8266 10600
rect 1104 10362 10028 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 10028 10362
rect 1104 10288 10028 10310
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3234 10248 3240 10260
rect 2731 10220 3240 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 4062 10248 4068 10260
rect 3651 10220 4068 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4985 10251 5043 10257
rect 4356 10220 4660 10248
rect 4356 10180 4384 10220
rect 3528 10152 4384 10180
rect 4632 10180 4660 10220
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5258 10248 5264 10260
rect 5031 10220 5264 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5810 10248 5816 10260
rect 5675 10220 5816 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 4893 10183 4951 10189
rect 4893 10180 4905 10183
rect 4632 10152 4905 10180
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 3326 10112 3332 10124
rect 3016 10084 3332 10112
rect 3016 10072 3022 10084
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 3528 10056 3556 10152
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 4356 10121 4384 10152
rect 4893 10149 4905 10152
rect 4939 10180 4951 10183
rect 5460 10180 5488 10211
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 6178 10248 6184 10260
rect 6135 10220 6184 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6638 10248 6644 10260
rect 6319 10220 6644 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6733 10251 6791 10257
rect 6733 10217 6745 10251
rect 6779 10248 6791 10251
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 6779 10220 7205 10248
rect 6779 10217 6791 10220
rect 6733 10211 6791 10217
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7193 10211 7251 10217
rect 7377 10251 7435 10257
rect 7377 10217 7389 10251
rect 7423 10248 7435 10251
rect 7558 10248 7564 10260
rect 7423 10220 7564 10248
rect 7423 10217 7435 10220
rect 7377 10211 7435 10217
rect 5721 10183 5779 10189
rect 5721 10180 5733 10183
rect 4939 10152 5733 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 5721 10149 5733 10152
rect 5767 10180 5779 10183
rect 6748 10180 6776 10211
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8021 10251 8079 10257
rect 8021 10248 8033 10251
rect 7800 10220 8033 10248
rect 7800 10208 7806 10220
rect 8021 10217 8033 10220
rect 8067 10217 8079 10251
rect 8021 10211 8079 10217
rect 5767 10152 6776 10180
rect 6917 10183 6975 10189
rect 5767 10149 5779 10152
rect 5721 10143 5779 10149
rect 6917 10149 6929 10183
rect 6963 10149 6975 10183
rect 6917 10143 6975 10149
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10081 4399 10115
rect 4341 10075 4399 10081
rect 4430 10072 4436 10124
rect 4488 10072 4494 10124
rect 4614 10072 4620 10124
rect 4672 10072 4678 10124
rect 6932 10112 6960 10143
rect 6932 10084 7512 10112
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3510 10044 3516 10056
rect 3467 10016 3516 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 2958 9936 2964 9988
rect 3016 9936 3022 9988
rect 3252 9976 3280 10007
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4856 10016 4997 10044
rect 4856 10004 4862 10016
rect 4985 10013 4997 10016
rect 5031 10044 5043 10047
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 5031 10016 5089 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 5077 10013 5089 10016
rect 5123 10044 5135 10047
rect 6178 10044 6184 10056
rect 5123 10016 6184 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 3602 9976 3608 9988
rect 3252 9948 3608 9976
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9945 4767 9979
rect 6380 9976 6408 10007
rect 7009 9979 7067 9985
rect 7009 9976 7021 9979
rect 4709 9939 4767 9945
rect 6104 9948 7021 9976
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 4246 9908 4252 9920
rect 3384 9880 4252 9908
rect 3384 9868 3390 9880
rect 4246 9868 4252 9880
rect 4304 9908 4310 9920
rect 4724 9908 4752 9939
rect 6104 9917 6132 9948
rect 7009 9945 7021 9948
rect 7055 9945 7067 9979
rect 7484 9976 7512 10084
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 7929 9979 7987 9985
rect 7929 9976 7941 9979
rect 7484 9948 7941 9976
rect 7009 9939 7067 9945
rect 7929 9945 7941 9948
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 4304 9880 5457 9908
rect 4304 9868 4310 9880
rect 5445 9877 5457 9880
rect 5491 9908 5503 9911
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 5491 9880 6101 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6089 9871 6147 9877
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6236 9880 6745 9908
rect 6236 9868 6242 9880
rect 6733 9877 6745 9880
rect 6779 9908 6791 9911
rect 7219 9911 7277 9917
rect 7219 9908 7231 9911
rect 6779 9880 7231 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 7219 9877 7231 9880
rect 7265 9908 7277 9911
rect 8220 9908 8248 10004
rect 7265 9880 8248 9908
rect 7265 9877 7277 9880
rect 7219 9871 7277 9877
rect 1104 9818 10028 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 10028 9818
rect 1104 9744 10028 9766
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 2096 9676 2912 9704
rect 2096 9664 2102 9676
rect 2884 9636 2912 9676
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3421 9707 3479 9713
rect 3421 9704 3433 9707
rect 3016 9676 3433 9704
rect 3016 9664 3022 9676
rect 3421 9673 3433 9676
rect 3467 9673 3479 9707
rect 3421 9667 3479 9673
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 4430 9704 4436 9716
rect 3660 9676 4436 9704
rect 3660 9664 3666 9676
rect 4430 9664 4436 9676
rect 4488 9704 4494 9716
rect 4798 9704 4804 9716
rect 4488 9676 4804 9704
rect 4488 9664 4494 9676
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 3510 9636 3516 9648
rect 2884 9608 3516 9636
rect 3510 9596 3516 9608
rect 3568 9636 3574 9648
rect 3568 9608 3832 9636
rect 3568 9596 3574 9608
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3804 9577 3832 9608
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3384 9540 3709 9568
rect 3384 9528 3390 9540
rect 3697 9537 3709 9540
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3602 9460 3608 9512
rect 3660 9460 3666 9512
rect 1104 9274 10028 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 10028 9274
rect 1104 9200 10028 9222
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 5902 9160 5908 9172
rect 4755 9132 5908 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 3237 9095 3295 9101
rect 3237 9092 3249 9095
rect 2740 9064 3249 9092
rect 2740 9052 2746 9064
rect 3237 9061 3249 9064
rect 3283 9061 3295 9095
rect 3237 9055 3295 9061
rect 5810 9024 5816 9036
rect 3436 8996 5816 9024
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 3436 8956 3464 8996
rect 5810 8984 5816 8996
rect 5868 9024 5874 9036
rect 5868 8996 8064 9024
rect 5868 8984 5874 8996
rect 1719 8928 3464 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1489 8891 1547 8897
rect 1489 8888 1501 8891
rect 992 8860 1501 8888
rect 992 8848 998 8860
rect 1489 8857 1501 8860
rect 1535 8857 1547 8891
rect 1489 8851 1547 8857
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8857 3295 8891
rect 3436 8888 3464 8928
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 5350 8956 5356 8968
rect 3559 8928 5356 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 6914 8956 6920 8968
rect 6687 8928 6920 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 8036 8900 8064 8996
rect 4157 8891 4215 8897
rect 4157 8888 4169 8891
rect 3436 8860 4169 8888
rect 3237 8851 3295 8857
rect 4157 8857 4169 8860
rect 4203 8857 4215 8891
rect 4157 8851 4215 8857
rect 4341 8891 4399 8897
rect 4341 8857 4353 8891
rect 4387 8888 4399 8891
rect 4430 8888 4436 8900
rect 4387 8860 4436 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 3252 8820 3280 8851
rect 4430 8848 4436 8860
rect 4488 8848 4494 8900
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 4614 8888 4620 8900
rect 4571 8860 4620 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 4724 8860 5290 8888
rect 3326 8820 3332 8832
rect 3252 8792 3332 8820
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3418 8780 3424 8832
rect 3476 8780 3482 8832
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 4028 8792 4077 8820
rect 4028 8780 4034 8792
rect 4065 8789 4077 8792
rect 4111 8820 4123 8823
rect 4724 8820 4752 8860
rect 8018 8848 8024 8900
rect 8076 8848 8082 8900
rect 4111 8792 4752 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4798 8780 4804 8832
rect 4856 8829 4862 8832
rect 4856 8823 4905 8829
rect 4856 8789 4859 8823
rect 4893 8789 4905 8823
rect 4856 8783 4905 8789
rect 4856 8780 4862 8783
rect 8662 8780 8668 8832
rect 8720 8829 8726 8832
rect 8720 8823 8769 8829
rect 8720 8789 8723 8823
rect 8757 8789 8769 8823
rect 8720 8783 8769 8789
rect 8720 8780 8726 8783
rect 1104 8730 10028 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 10028 8730
rect 1104 8656 10028 8678
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 5162 8619 5220 8625
rect 3476 8588 5120 8616
rect 3476 8576 3482 8588
rect 3970 8548 3976 8560
rect 3726 8520 3976 8548
rect 3970 8508 3976 8520
rect 4028 8508 4034 8560
rect 2682 8440 2688 8492
rect 2740 8440 2746 8492
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4798 8480 4804 8492
rect 4571 8452 4804 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5092 8489 5120 8588
rect 5162 8585 5174 8619
rect 5208 8616 5220 8619
rect 6270 8616 6276 8628
rect 5208 8588 6276 8616
rect 5208 8585 5220 8588
rect 5162 8579 5220 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6564 8588 7236 8616
rect 5276 8520 6500 8548
rect 5276 8489 5304 8520
rect 6472 8492 6500 8520
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 2314 8372 2320 8424
rect 2372 8372 2378 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8381 4675 8415
rect 4617 8375 4675 8381
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8412 4951 8415
rect 5000 8412 5028 8443
rect 4939 8384 5028 8412
rect 4939 8381 4951 8384
rect 4893 8375 4951 8381
rect 4632 8344 4660 8375
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 5368 8412 5396 8443
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5500 8452 5549 8480
rect 5500 8440 5506 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5806 8483 5864 8489
rect 5806 8449 5818 8483
rect 5852 8449 5864 8483
rect 5806 8443 5864 8449
rect 5644 8412 5672 8443
rect 5224 8384 5396 8412
rect 5460 8384 5672 8412
rect 5828 8412 5856 8443
rect 6454 8440 6460 8492
rect 6512 8440 6518 8492
rect 6564 8480 6592 8588
rect 7208 8557 7236 8588
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 8849 8619 8907 8625
rect 8849 8616 8861 8619
rect 7340 8588 8861 8616
rect 7340 8576 7346 8588
rect 8849 8585 8861 8588
rect 8895 8585 8907 8619
rect 8849 8579 8907 8585
rect 6641 8551 6699 8557
rect 6641 8517 6653 8551
rect 6687 8548 6699 8551
rect 7193 8551 7251 8557
rect 6687 8520 7144 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6564 8452 6745 8480
rect 6733 8449 6745 8452
rect 6779 8480 6791 8483
rect 6822 8480 6828 8492
rect 6779 8452 6828 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7116 8480 7144 8520
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 7239 8520 8524 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 7944 8489 7972 8520
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7116 8452 7849 8480
rect 7300 8424 7328 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 5902 8412 5908 8424
rect 5828 8384 5908 8412
rect 5224 8372 5230 8384
rect 5460 8353 5488 8384
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 7282 8372 7288 8424
rect 7340 8372 7346 8424
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 5445 8347 5503 8353
rect 5445 8344 5457 8347
rect 4632 8316 5457 8344
rect 5445 8313 5457 8316
rect 5491 8313 5503 8347
rect 5445 8307 5503 8313
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 7006 8344 7012 8356
rect 6871 8316 7012 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 7006 8304 7012 8316
rect 7064 8344 7070 8356
rect 7484 8344 7512 8375
rect 7064 8316 7512 8344
rect 7064 8304 7070 8316
rect 4111 8279 4169 8285
rect 4111 8245 4123 8279
rect 4157 8276 4169 8279
rect 4706 8276 4712 8288
rect 4157 8248 4712 8276
rect 4157 8245 4169 8248
rect 4111 8239 4169 8245
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 5408 8248 5733 8276
rect 5408 8236 5414 8248
rect 5721 8245 5733 8248
rect 5767 8245 5779 8279
rect 5721 8239 5779 8245
rect 6457 8279 6515 8285
rect 6457 8245 6469 8279
rect 6503 8276 6515 8279
rect 7098 8276 7104 8288
rect 6503 8248 7104 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 7193 8279 7251 8285
rect 7193 8245 7205 8279
rect 7239 8276 7251 8279
rect 7282 8276 7288 8288
rect 7239 8248 7288 8276
rect 7239 8245 7251 8248
rect 7193 8239 7251 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 7374 8236 7380 8288
rect 7432 8236 7438 8288
rect 7650 8236 7656 8288
rect 7708 8236 7714 8288
rect 8404 8276 8432 8443
rect 8496 8421 8524 8520
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9364 8452 9413 8480
rect 9364 8440 9370 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 9232 8412 9260 8440
rect 8527 8384 9260 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 8803 8316 9229 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 9217 8307 9275 8313
rect 9582 8304 9588 8356
rect 9640 8304 9646 8356
rect 8662 8276 8668 8288
rect 8404 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8276 8726 8288
rect 9306 8276 9312 8288
rect 8720 8248 9312 8276
rect 8720 8236 8726 8248
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 1104 8186 10028 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 10028 8186
rect 1104 8112 10028 8134
rect 5399 8075 5457 8081
rect 5399 8041 5411 8075
rect 5445 8072 5457 8075
rect 7006 8072 7012 8084
rect 5445 8044 7012 8072
rect 5445 8041 5457 8044
rect 5399 8035 5457 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 8202 8072 8208 8084
rect 8036 8044 8208 8072
rect 4706 7964 4712 8016
rect 4764 8004 4770 8016
rect 5261 8007 5319 8013
rect 5261 8004 5273 8007
rect 4764 7976 5273 8004
rect 4764 7964 4770 7976
rect 5261 7973 5273 7976
rect 5307 7973 5319 8007
rect 5261 7967 5319 7973
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2314 7936 2320 7948
rect 1811 7908 2320 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2314 7896 2320 7908
rect 2372 7936 2378 7948
rect 3694 7936 3700 7948
rect 2372 7908 3700 7936
rect 2372 7896 2378 7908
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4614 7936 4620 7948
rect 4479 7908 4620 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 2130 7828 2136 7880
rect 2188 7828 2194 7880
rect 3559 7871 3617 7877
rect 3559 7837 3571 7871
rect 3605 7868 3617 7871
rect 4154 7868 4160 7880
rect 3605 7840 4160 7868
rect 3605 7837 3617 7840
rect 3559 7831 3617 7837
rect 4154 7828 4160 7840
rect 4212 7868 4218 7880
rect 4448 7868 4476 7899
rect 4614 7896 4620 7908
rect 4672 7936 4678 7948
rect 5166 7936 5172 7948
rect 4672 7908 5172 7936
rect 4672 7896 4678 7908
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5276 7936 5304 7967
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7561 8007 7619 8013
rect 7561 8004 7573 8007
rect 7432 7976 7573 8004
rect 7432 7964 7438 7976
rect 7561 7973 7573 7976
rect 7607 7973 7619 8007
rect 7561 7967 7619 7973
rect 7650 7964 7656 8016
rect 7708 7964 7714 8016
rect 8036 8004 8064 8044
rect 8202 8032 8208 8044
rect 8260 8072 8266 8084
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8260 8044 8677 8072
rect 8260 8032 8266 8044
rect 8665 8041 8677 8044
rect 8711 8072 8723 8075
rect 9030 8072 9036 8084
rect 8711 8044 9036 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 7760 7976 8064 8004
rect 5442 7936 5448 7948
rect 5276 7908 5448 7936
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7190 7936 7196 7948
rect 6972 7908 7196 7936
rect 6972 7896 6978 7908
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 4212 7840 4476 7868
rect 4985 7871 5043 7877
rect 4212 7828 4218 7840
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5350 7868 5356 7880
rect 5031 7840 5356 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 6871 7840 7297 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 7760 7877 7788 7976
rect 8110 7964 8116 8016
rect 8168 8004 8174 8016
rect 9493 8007 9551 8013
rect 9493 8004 9505 8007
rect 8168 7976 9505 8004
rect 8168 7964 8174 7976
rect 9493 7973 9505 7976
rect 9539 7973 9551 8007
rect 9493 7967 9551 7973
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8128 7908 8953 7936
rect 8128 7877 8156 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8343 7871 8401 7877
rect 8343 7837 8355 7871
rect 8389 7868 8401 7871
rect 8478 7868 8484 7880
rect 8389 7840 8484 7868
rect 8389 7837 8401 7840
rect 8343 7831 8401 7837
rect 3970 7800 3976 7812
rect 3174 7772 3976 7800
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 4709 7803 4767 7809
rect 4709 7769 4721 7803
rect 4755 7800 4767 7803
rect 5442 7800 5448 7812
rect 4755 7772 5448 7800
rect 4755 7769 4767 7772
rect 4709 7763 4767 7769
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 5810 7760 5816 7812
rect 5868 7760 5874 7812
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7944 7800 7972 7831
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9272 7840 9413 7868
rect 9272 7828 9278 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9723 7840 10180 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 7156 7772 7972 7800
rect 7156 7760 7162 7772
rect 8202 7760 8208 7812
rect 8260 7760 8266 7812
rect 10152 7744 10180 7840
rect 3786 7692 3792 7744
rect 3844 7692 3850 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 4893 7735 4951 7741
rect 4893 7732 4905 7735
rect 4856 7704 4905 7732
rect 4856 7692 4862 7704
rect 4893 7701 4905 7704
rect 4939 7701 4951 7735
rect 4893 7695 4951 7701
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 5166 7732 5172 7744
rect 5123 7704 5172 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 8352 7704 8493 7732
rect 8352 7692 8358 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 9306 7692 9312 7744
rect 9364 7692 9370 7744
rect 10134 7692 10140 7744
rect 10192 7692 10198 7744
rect 1104 7642 10028 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 10028 7642
rect 1104 7568 10028 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 3145 7531 3203 7537
rect 2188 7500 2774 7528
rect 2188 7488 2194 7500
rect 2746 7256 2774 7500
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3786 7528 3792 7540
rect 3191 7500 3792 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 3970 7488 3976 7540
rect 4028 7528 4034 7540
rect 6457 7531 6515 7537
rect 4028 7500 4384 7528
rect 4028 7488 4034 7500
rect 3418 7460 3424 7472
rect 3252 7432 3424 7460
rect 3252 7401 3280 7432
rect 3418 7420 3424 7432
rect 3476 7460 3482 7472
rect 3513 7463 3571 7469
rect 3513 7460 3525 7463
rect 3476 7432 3525 7460
rect 3476 7420 3482 7432
rect 3513 7429 3525 7432
rect 3559 7429 3571 7463
rect 4356 7460 4384 7500
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 6638 7528 6644 7540
rect 6503 7500 6644 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 7064 7500 7113 7528
rect 7064 7488 7070 7500
rect 7101 7497 7113 7500
rect 7147 7497 7159 7531
rect 7101 7491 7159 7497
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 8938 7528 8944 7540
rect 7340 7500 8944 7528
rect 7340 7488 7346 7500
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9631 7531 9689 7537
rect 9631 7528 9643 7531
rect 9180 7500 9643 7528
rect 9180 7488 9186 7500
rect 9631 7497 9643 7500
rect 9677 7497 9689 7531
rect 9631 7491 9689 7497
rect 6914 7460 6920 7472
rect 3513 7423 3571 7429
rect 3620 7432 3832 7460
rect 4356 7432 4462 7460
rect 6656 7432 6920 7460
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 2976 7324 3004 7355
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 3620 7401 3648 7432
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3694 7352 3700 7404
rect 3752 7352 3758 7404
rect 3804 7392 3832 7432
rect 6365 7395 6423 7401
rect 3804 7364 4200 7392
rect 3344 7324 3372 7352
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 2976 7296 3372 7324
rect 3712 7296 4077 7324
rect 2961 7259 3019 7265
rect 2961 7256 2973 7259
rect 2746 7228 2973 7256
rect 2961 7225 2973 7228
rect 3007 7225 3019 7259
rect 2961 7219 3019 7225
rect 3329 7259 3387 7265
rect 3329 7225 3341 7259
rect 3375 7256 3387 7259
rect 3712 7256 3740 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4172 7324 4200 7364
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6546 7392 6552 7404
rect 6411 7364 6552 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 6656 7401 6684 7432
rect 6914 7420 6920 7432
rect 6972 7460 6978 7472
rect 6972 7432 7328 7460
rect 6972 7420 6978 7432
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7300 7392 7328 7432
rect 7466 7420 7472 7472
rect 7524 7420 7530 7472
rect 8110 7392 8116 7404
rect 7300 7364 8116 7392
rect 7193 7355 7251 7361
rect 5258 7324 5264 7336
rect 4172 7296 5264 7324
rect 4065 7287 4123 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 6564 7324 6592 7352
rect 7208 7324 7236 7355
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8294 7392 8300 7404
rect 8251 7364 8300 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 7834 7324 7840 7336
rect 6564 7296 7236 7324
rect 7760 7296 7840 7324
rect 3375 7228 3740 7256
rect 3375 7225 3387 7228
rect 3329 7219 3387 7225
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 6917 7259 6975 7265
rect 6917 7256 6929 7259
rect 6696 7228 6929 7256
rect 6696 7216 6702 7228
rect 6917 7225 6929 7228
rect 6963 7225 6975 7259
rect 6917 7219 6975 7225
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 7760 7256 7788 7296
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8956 7324 8984 7446
rect 8076 7296 8984 7324
rect 8076 7284 8082 7296
rect 7248 7228 7788 7256
rect 7248 7216 7254 7228
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5350 7188 5356 7200
rect 4948 7160 5356 7188
rect 4948 7148 4954 7160
rect 5350 7148 5356 7160
rect 5408 7188 5414 7200
rect 5491 7191 5549 7197
rect 5491 7188 5503 7191
rect 5408 7160 5503 7188
rect 5408 7148 5414 7160
rect 5491 7157 5503 7160
rect 5537 7157 5549 7191
rect 5491 7151 5549 7157
rect 1104 7098 10028 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 10028 7098
rect 1104 7024 10028 7046
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 8294 6984 8300 6996
rect 7892 6956 8300 6984
rect 7892 6944 7898 6956
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8938 6944 8944 6996
rect 8996 6944 9002 6996
rect 4890 6916 4896 6928
rect 4172 6888 4896 6916
rect 4172 6857 4200 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4338 6808 4344 6860
rect 4396 6808 4402 6860
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4798 6848 4804 6860
rect 4479 6820 4804 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 9306 6808 9312 6860
rect 9364 6808 9370 6860
rect 3418 6740 3424 6792
rect 3476 6780 3482 6792
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3476 6752 3525 6780
rect 3476 6740 3482 6752
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3602 6740 3608 6792
rect 3660 6740 3666 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 4062 6712 4068 6724
rect 3384 6684 4068 6712
rect 3384 6672 3390 6684
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 4264 6712 4292 6743
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4672 6752 5089 6780
rect 4672 6740 4678 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 6454 6740 6460 6792
rect 6512 6780 6518 6792
rect 7650 6780 7656 6792
rect 6512 6752 7656 6780
rect 6512 6740 6518 6752
rect 7650 6740 7656 6752
rect 7708 6780 7714 6792
rect 8570 6780 8576 6792
rect 7708 6752 8576 6780
rect 7708 6740 7714 6752
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 4706 6712 4712 6724
rect 4264 6684 4712 6712
rect 4706 6672 4712 6684
rect 4764 6672 4770 6724
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6380 6684 7021 6712
rect 6380 6656 6408 6684
rect 7009 6681 7021 6684
rect 7055 6681 7067 6715
rect 7009 6675 7067 6681
rect 3418 6604 3424 6656
rect 3476 6653 3482 6656
rect 3476 6607 3485 6653
rect 3476 6604 3482 6607
rect 4614 6604 4620 6656
rect 4672 6604 4678 6656
rect 6362 6604 6368 6656
rect 6420 6604 6426 6656
rect 9582 6604 9588 6656
rect 9640 6604 9646 6656
rect 1104 6554 10028 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 10028 6554
rect 1104 6480 10028 6502
rect 3694 6440 3700 6452
rect 3068 6412 3700 6440
rect 3068 6316 3096 6412
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 4614 6400 4620 6452
rect 4672 6400 4678 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5258 6440 5264 6452
rect 5031 6412 5264 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 6454 6440 6460 6452
rect 5684 6412 6460 6440
rect 5684 6400 5690 6412
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 8478 6400 8484 6452
rect 8536 6400 8542 6452
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 4632 6304 4660 6400
rect 4798 6332 4804 6384
rect 4856 6381 4862 6384
rect 4856 6375 4905 6381
rect 4856 6341 4859 6375
rect 4893 6372 4905 6375
rect 8496 6372 8524 6400
rect 4893 6344 6040 6372
rect 4893 6341 4905 6344
rect 4856 6335 4905 6341
rect 4856 6332 4862 6335
rect 5199 6307 5257 6313
rect 5199 6304 5211 6307
rect 4632 6276 5211 6304
rect 5199 6273 5211 6276
rect 5245 6273 5257 6307
rect 5199 6267 5257 6273
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 5074 6236 5080 6248
rect 4672 6208 5080 6236
rect 4672 6196 4678 6208
rect 5074 6196 5080 6208
rect 5132 6236 5138 6248
rect 5368 6236 5396 6264
rect 5132 6208 5396 6236
rect 5132 6196 5138 6208
rect 5460 6112 5488 6267
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6012 6313 6040 6344
rect 7300 6344 9076 6372
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5592 6276 5825 6304
rect 5592 6264 5598 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 6638 6304 6644 6316
rect 6595 6276 6644 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7300 6313 7328 6344
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6972 6276 7021 6304
rect 6972 6264 6978 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 6454 6196 6460 6248
rect 6512 6196 6518 6248
rect 8478 6196 8484 6248
rect 8536 6196 8542 6248
rect 8938 6196 8944 6248
rect 8996 6196 9002 6248
rect 6914 6128 6920 6180
rect 6972 6128 6978 6180
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 7374 6168 7380 6180
rect 7331 6140 7380 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 8496 6168 8524 6196
rect 9048 6180 9076 6344
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 9692 6236 9720 6267
rect 10134 6236 10140 6248
rect 9692 6208 10140 6236
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 8496 6140 8984 6168
rect 2222 6060 2228 6112
rect 2280 6060 2286 6112
rect 5442 6060 5448 6112
rect 5500 6060 5506 6112
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 8846 6060 8852 6112
rect 8904 6060 8910 6112
rect 8956 6100 8984 6140
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9217 6171 9275 6177
rect 9217 6168 9229 6171
rect 9088 6140 9229 6168
rect 9088 6128 9094 6140
rect 9217 6137 9229 6140
rect 9263 6137 9275 6171
rect 9217 6131 9275 6137
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 8956 6072 9505 6100
rect 9493 6069 9505 6072
rect 9539 6069 9551 6103
rect 9493 6063 9551 6069
rect 1104 6010 10028 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 10028 6010
rect 1104 5936 10028 5958
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3660 5868 3893 5896
rect 3660 5856 3666 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4706 5896 4712 5908
rect 4387 5868 4712 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4356 5828 4384 5859
rect 4706 5856 4712 5868
rect 4764 5896 4770 5908
rect 5353 5899 5411 5905
rect 4764 5868 4936 5896
rect 4764 5856 4770 5868
rect 4080 5800 4384 5828
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 3050 5760 3056 5772
rect 1811 5732 3056 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2222 5692 2228 5704
rect 2179 5664 2228 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 4080 5701 4108 5800
rect 4798 5788 4804 5840
rect 4856 5788 4862 5840
rect 4908 5828 4936 5868
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 6454 5896 6460 5908
rect 5399 5868 6460 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 6638 5856 6644 5908
rect 6696 5905 6702 5908
rect 6696 5899 6745 5905
rect 6696 5865 6699 5899
rect 6733 5865 6745 5899
rect 6696 5859 6745 5865
rect 6696 5856 6702 5859
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8536 5868 9045 5896
rect 8536 5856 8542 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 4908 5800 6592 5828
rect 5810 5760 5816 5772
rect 4264 5732 5816 5760
rect 4264 5701 4292 5732
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5760 6147 5763
rect 6135 5732 6500 5760
rect 6135 5729 6147 5732
rect 6089 5723 6147 5729
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4614 5692 4620 5704
rect 4571 5664 4620 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4798 5692 4804 5704
rect 4755 5664 4804 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5442 5692 5448 5704
rect 4908 5664 5448 5692
rect 2866 5584 2872 5636
rect 2924 5584 2930 5636
rect 4264 5596 4752 5624
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 3559 5559 3617 5565
rect 3559 5525 3571 5559
rect 3605 5556 3617 5559
rect 4264 5556 4292 5596
rect 3605 5528 4292 5556
rect 4724 5556 4752 5596
rect 4908 5556 4936 5664
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 5074 5584 5080 5636
rect 5132 5584 5138 5636
rect 5169 5627 5227 5633
rect 5169 5593 5181 5627
rect 5215 5624 5227 5627
rect 6178 5624 6184 5636
rect 5215 5596 6184 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 6178 5584 6184 5596
rect 6236 5624 6242 5636
rect 6380 5624 6408 5655
rect 6236 5596 6408 5624
rect 6472 5624 6500 5732
rect 6564 5701 6592 5800
rect 8938 5788 8944 5840
rect 8996 5788 9002 5840
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8352 5732 8493 5760
rect 8352 5720 8358 5732
rect 8481 5729 8493 5732
rect 8527 5729 8539 5763
rect 8956 5760 8984 5788
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 8956 5732 9229 5760
rect 8481 5723 8539 5729
rect 9217 5729 9229 5732
rect 9263 5760 9275 5763
rect 9674 5760 9680 5772
rect 9263 5732 9680 5760
rect 9263 5729 9275 5732
rect 9217 5723 9275 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9030 5692 9036 5704
rect 8987 5664 9036 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 8588 5624 8616 5655
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9582 5624 9588 5636
rect 6472 5596 7052 5624
rect 7774 5596 7880 5624
rect 8588 5596 9588 5624
rect 6236 5584 6242 5596
rect 4724 5528 4936 5556
rect 4985 5559 5043 5565
rect 3605 5525 3617 5528
rect 3559 5519 3617 5525
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 6270 5556 6276 5568
rect 5031 5528 6276 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6454 5516 6460 5568
rect 6512 5516 6518 5568
rect 7024 5556 7052 5596
rect 7190 5556 7196 5568
rect 7024 5528 7196 5556
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 7852 5556 7880 5596
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 8018 5556 8024 5568
rect 7852 5528 8024 5556
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8754 5516 8760 5568
rect 8812 5516 8818 5568
rect 9490 5516 9496 5568
rect 9548 5516 9554 5568
rect 1104 5466 10028 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 10028 5466
rect 1104 5392 10028 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 2866 5352 2872 5364
rect 2823 5324 2872 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 3108 5324 3157 5352
rect 3108 5312 3114 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 3145 5315 3203 5321
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 3568 5324 4997 5352
rect 3568 5312 3574 5324
rect 4985 5321 4997 5324
rect 5031 5352 5043 5355
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 5031 5324 7113 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 7101 5321 7113 5324
rect 7147 5352 7159 5355
rect 7374 5352 7380 5364
rect 7147 5324 7380 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7374 5312 7380 5324
rect 7432 5352 7438 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 7432 5324 7481 5352
rect 7432 5312 7438 5324
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 7469 5315 7527 5321
rect 8110 5312 8116 5364
rect 8168 5312 8174 5364
rect 9674 5312 9680 5364
rect 9732 5312 9738 5364
rect 4617 5287 4675 5293
rect 4617 5253 4629 5287
rect 4663 5284 4675 5287
rect 6362 5284 6368 5296
rect 4663 5256 6368 5284
rect 4663 5253 4675 5256
rect 4617 5247 4675 5253
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 7248 5256 7297 5284
rect 7248 5244 7254 5256
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 7285 5247 7343 5253
rect 7650 5244 7656 5296
rect 7708 5244 7714 5296
rect 8128 5284 8156 5312
rect 7760 5256 8156 5284
rect 8205 5287 8263 5293
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 4062 5216 4068 5228
rect 3384 5188 4068 5216
rect 3384 5176 3390 5188
rect 4062 5176 4068 5188
rect 4120 5216 4126 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4120 5188 4813 5216
rect 4120 5176 4126 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 2130 5108 2136 5160
rect 2188 5108 2194 5160
rect 4816 5080 4844 5179
rect 5092 5148 5120 5179
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5675 5188 6009 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 5997 5185 6009 5188
rect 6043 5216 6055 5219
rect 6043 5188 6132 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 5258 5148 5264 5160
rect 5092 5120 5264 5148
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5552 5148 5580 5176
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5552 5120 5825 5148
rect 5813 5117 5825 5120
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 5626 5080 5632 5092
rect 4816 5052 5632 5080
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 6104 5024 6132 5188
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6328 5188 6561 5216
rect 6328 5176 6334 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6932 5216 6960 5244
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6932 5188 7021 5216
rect 6549 5179 6607 5185
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 6454 5108 6460 5160
rect 6512 5108 6518 5160
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 7392 5148 7420 5179
rect 6963 5120 7420 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 7285 5083 7343 5089
rect 7285 5049 7297 5083
rect 7331 5080 7343 5083
rect 7760 5080 7788 5256
rect 8205 5253 8217 5287
rect 8251 5284 8263 5287
rect 8478 5284 8484 5296
rect 8251 5256 8484 5284
rect 8251 5253 8263 5256
rect 8205 5247 8263 5253
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 8846 5244 8852 5296
rect 8904 5244 8910 5296
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8294 5148 8300 5160
rect 7975 5120 8300 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 7331 5052 7788 5080
rect 7331 5049 7343 5052
rect 7285 5043 7343 5049
rect 4801 5015 4859 5021
rect 4801 4981 4813 5015
rect 4847 5012 4859 5015
rect 4982 5012 4988 5024
rect 4847 4984 4988 5012
rect 4847 4981 4859 4984
rect 4801 4975 4859 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5169 5015 5227 5021
rect 5169 4981 5181 5015
rect 5215 5012 5227 5015
rect 5258 5012 5264 5024
rect 5215 4984 5264 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6086 4972 6092 5024
rect 6144 4972 6150 5024
rect 7653 5015 7711 5021
rect 7653 4981 7665 5015
rect 7699 5012 7711 5015
rect 8202 5012 8208 5024
rect 7699 4984 8208 5012
rect 7699 4981 7711 4984
rect 7653 4975 7711 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 1104 4922 10028 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 10028 4922
rect 1104 4848 10028 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 2130 4808 2136 4820
rect 1443 4780 2136 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 3050 4768 3056 4820
rect 3108 4768 3114 4820
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 5442 4808 5448 4820
rect 4948 4780 5448 4808
rect 4948 4768 4954 4780
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6503 4811 6561 4817
rect 6503 4808 6515 4811
rect 6144 4780 6515 4808
rect 6144 4768 6150 4780
rect 6503 4777 6515 4780
rect 6549 4777 6561 4811
rect 6503 4771 6561 4777
rect 3068 4672 3096 4768
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3418 4740 3424 4752
rect 3375 4712 3424 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 3418 4700 3424 4712
rect 3476 4700 3482 4752
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6779 4743 6837 4749
rect 6779 4740 6791 4743
rect 6328 4712 6791 4740
rect 6328 4700 6334 4712
rect 6779 4709 6791 4712
rect 6825 4709 6837 4743
rect 6779 4703 6837 4709
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 3068 4644 3157 4672
rect 3145 4641 3157 4644
rect 3191 4672 3203 4675
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 3191 4644 4721 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 4709 4641 4721 4644
rect 4755 4641 4767 4675
rect 4709 4635 4767 4641
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5077 4675 5135 4681
rect 5077 4672 5089 4675
rect 5040 4644 5089 4672
rect 5040 4632 5046 4644
rect 5077 4641 5089 4644
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8573 4675 8631 4681
rect 8573 4672 8585 4675
rect 8352 4644 8585 4672
rect 8352 4632 8358 4644
rect 8573 4641 8585 4644
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8812 4644 9045 4672
rect 8812 4632 8818 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4672 9367 4675
rect 9490 4672 9496 4684
rect 9355 4644 9496 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 3326 4564 3332 4616
rect 3384 4564 3390 4616
rect 3510 4564 3516 4616
rect 3568 4564 3574 4616
rect 3602 4564 3608 4616
rect 3660 4564 3666 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4614 4604 4620 4616
rect 4479 4576 4620 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 8202 4564 8208 4616
rect 8260 4564 8266 4616
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 2130 4496 2136 4548
rect 2188 4496 2194 4548
rect 2869 4539 2927 4545
rect 2869 4505 2881 4539
rect 2915 4505 2927 4539
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 2869 4499 2927 4505
rect 3436 4508 3801 4536
rect 2884 4468 2912 4499
rect 3436 4468 3464 4508
rect 3789 4505 3801 4508
rect 3835 4505 3847 4539
rect 6118 4508 6224 4536
rect 7866 4508 7972 4536
rect 3789 4499 3847 4505
rect 2884 4440 3464 4468
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 4798 4468 4804 4480
rect 4028 4440 4804 4468
rect 4028 4428 4034 4440
rect 4798 4428 4804 4440
rect 4856 4468 4862 4480
rect 6196 4468 6224 4508
rect 7944 4468 7972 4508
rect 8662 4468 8668 4480
rect 4856 4440 8668 4468
rect 4856 4428 4862 4440
rect 8662 4428 8668 4440
rect 8720 4468 8726 4480
rect 9140 4468 9168 4567
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 8720 4440 9168 4468
rect 8720 4428 8726 4440
rect 9490 4428 9496 4480
rect 9548 4428 9554 4480
rect 1104 4378 10028 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 10028 4378
rect 1104 4304 10028 4326
rect 2130 4224 2136 4276
rect 2188 4224 2194 4276
rect 4798 4224 4804 4276
rect 4856 4224 4862 4276
rect 5258 4224 5264 4276
rect 5316 4224 5322 4276
rect 5350 4224 5356 4276
rect 5408 4224 5414 4276
rect 9214 4224 9220 4276
rect 9272 4224 9278 4276
rect 4816 4196 4844 4224
rect 4554 4168 4844 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 2225 4131 2283 4137
rect 2225 4128 2237 4131
rect 1596 4100 2237 4128
rect 1596 4001 1624 4100
rect 2225 4097 2237 4100
rect 2271 4128 2283 4131
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 2271 4100 2329 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 3108 4100 3157 4128
rect 3108 4088 3114 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 5276 4137 5304 4224
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 3476 4100 3525 4128
rect 3476 4088 3482 4100
rect 3513 4097 3525 4100
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 6454 4128 6460 4140
rect 5491 4100 6460 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 9048 4100 9137 4128
rect 4939 4063 4997 4069
rect 4939 4029 4951 4063
rect 4985 4060 4997 4063
rect 5534 4060 5540 4072
rect 4985 4032 5540 4060
rect 4985 4029 4997 4032
rect 4939 4023 4997 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 9048 4001 9076 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9490 4128 9496 4140
rect 9447 4100 9496 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3961 1639 3995
rect 1581 3955 1639 3961
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 2406 3884 2412 3936
rect 2464 3884 2470 3936
rect 9582 3884 9588 3936
rect 9640 3884 9646 3936
rect 1104 3834 10028 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 10028 3834
rect 1104 3760 10028 3782
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3660 3692 4077 3720
rect 3660 3680 3666 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4614 3680 4620 3732
rect 4672 3680 4678 3732
rect 3145 3655 3203 3661
rect 3145 3621 3157 3655
rect 3191 3652 3203 3655
rect 4632 3652 4660 3680
rect 3191 3624 4660 3652
rect 3191 3621 3203 3624
rect 3145 3615 3203 3621
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 3050 3584 3056 3596
rect 1443 3556 3056 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 4706 3584 4712 3596
rect 4479 3556 4712 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 5534 3516 5540 3528
rect 4387 3488 5540 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 7883 3488 7972 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 1578 3408 1584 3460
rect 1636 3448 1642 3460
rect 1673 3451 1731 3457
rect 1673 3448 1685 3451
rect 1636 3420 1685 3448
rect 1636 3408 1642 3420
rect 1673 3417 1685 3420
rect 1719 3417 1731 3451
rect 1673 3411 1731 3417
rect 2406 3408 2412 3460
rect 2464 3408 2470 3460
rect 7558 3408 7564 3460
rect 7616 3408 7622 3460
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 7760 3380 7788 3479
rect 7944 3392 7972 3488
rect 7524 3352 7788 3380
rect 7524 3340 7530 3352
rect 7834 3340 7840 3392
rect 7892 3340 7898 3392
rect 7926 3340 7932 3392
rect 7984 3340 7990 3392
rect 1104 3290 10028 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 10028 3290
rect 1104 3216 10028 3238
rect 7558 3176 7564 3188
rect 6932 3148 7564 3176
rect 6638 3108 6644 3120
rect 5920 3080 6644 3108
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4798 3040 4804 3052
rect 4479 3012 4804 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 4982 3000 4988 3052
rect 5040 3000 5046 3052
rect 5920 3040 5948 3080
rect 6638 3068 6644 3080
rect 6696 3108 6702 3120
rect 6932 3117 6960 3148
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 7892 3148 9444 3176
rect 7892 3136 7898 3148
rect 6917 3111 6975 3117
rect 6917 3108 6929 3111
rect 6696 3080 6929 3108
rect 6696 3068 6702 3080
rect 6917 3077 6929 3080
rect 6963 3077 6975 3111
rect 6917 3071 6975 3077
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 7926 3108 7932 3120
rect 7248 3080 7932 3108
rect 7248 3068 7254 3080
rect 7926 3068 7932 3080
rect 7984 3108 7990 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7984 3080 8217 3108
rect 7984 3068 7990 3080
rect 8205 3077 8217 3080
rect 8251 3108 8263 3111
rect 8633 3111 8691 3117
rect 8633 3108 8645 3111
rect 8251 3080 8645 3108
rect 8251 3077 8263 3080
rect 8205 3071 8263 3077
rect 8633 3077 8645 3080
rect 8679 3077 8691 3111
rect 8633 3071 8691 3077
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3077 8907 3111
rect 8849 3071 8907 3077
rect 5828 3012 5948 3040
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 5828 2981 5856 3012
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6104 3012 6561 3040
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4212 2944 4261 2972
rect 4212 2932 4218 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2972 4399 2975
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4387 2944 4905 2972
rect 4387 2941 4399 2944
rect 4341 2935 4399 2941
rect 4893 2941 4905 2944
rect 4939 2972 4951 2975
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 4939 2944 5825 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5813 2941 5825 2944
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 5905 2975 5963 2981
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 6104 2972 6132 3012
rect 6549 3009 6561 3012
rect 6595 3040 6607 3043
rect 7466 3040 7472 3052
rect 6595 3012 7472 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7616 3012 7849 3040
rect 7616 3000 7622 3012
rect 7837 3009 7849 3012
rect 7883 3040 7895 3043
rect 8864 3040 8892 3071
rect 9416 3049 9444 3148
rect 7883 3012 8892 3040
rect 9401 3043 9459 3049
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 5951 2944 6132 2972
rect 6181 2975 6239 2981
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 7098 2972 7104 2984
rect 6227 2944 7104 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 4264 2904 4292 2935
rect 4982 2904 4988 2916
rect 4264 2876 4988 2904
rect 4982 2864 4988 2876
rect 5040 2904 5046 2916
rect 5920 2904 5948 2935
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7190 2904 7196 2916
rect 5040 2876 5948 2904
rect 6932 2876 7196 2904
rect 5040 2864 5046 2876
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 3752 2808 4077 2836
rect 3752 2796 3758 2808
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4065 2799 4123 2805
rect 4614 2796 4620 2848
rect 4672 2796 4678 2848
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 6932 2845 6960 2876
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 7484 2904 7512 3000
rect 7484 2876 8708 2904
rect 6917 2839 6975 2845
rect 6917 2836 6929 2839
rect 6052 2808 6929 2836
rect 6052 2796 6058 2808
rect 6917 2805 6929 2808
rect 6963 2805 6975 2839
rect 6917 2799 6975 2805
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 7374 2836 7380 2848
rect 7147 2808 7380 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7484 2836 7512 2876
rect 7561 2839 7619 2845
rect 7561 2836 7573 2839
rect 7484 2808 7573 2836
rect 7561 2805 7573 2808
rect 7607 2805 7619 2839
rect 7561 2799 7619 2805
rect 7742 2796 7748 2848
rect 7800 2796 7806 2848
rect 8220 2845 8248 2876
rect 8205 2839 8263 2845
rect 8205 2805 8217 2839
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 8386 2796 8392 2848
rect 8444 2796 8450 2848
rect 8478 2796 8484 2848
rect 8536 2796 8542 2848
rect 8680 2845 8708 2876
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 9585 2839 9643 2845
rect 9585 2805 9597 2839
rect 9631 2836 9643 2839
rect 9674 2836 9680 2848
rect 9631 2808 9680 2836
rect 9631 2805 9643 2808
rect 9585 2799 9643 2805
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 1104 2746 10028 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 10028 2746
rect 1104 2672 10028 2694
rect 4798 2592 4804 2644
rect 4856 2592 4862 2644
rect 6638 2592 6644 2644
rect 6696 2592 6702 2644
rect 4062 2456 4068 2508
rect 4120 2456 4126 2508
rect 4816 2496 4844 2592
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 4816 2468 5549 2496
rect 5537 2465 5549 2468
rect 5583 2496 5595 2499
rect 5994 2496 6000 2508
rect 5583 2468 6000 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6656 2505 6684 2592
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 7837 2567 7895 2573
rect 7837 2564 7849 2567
rect 7156 2536 7849 2564
rect 7156 2524 7162 2536
rect 7837 2533 7849 2536
rect 7883 2533 7895 2567
rect 7837 2527 7895 2533
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2465 6699 2499
rect 6641 2459 6699 2465
rect 8404 2468 9168 2496
rect 8404 2440 8432 2468
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3694 2428 3700 2440
rect 3651 2400 3700 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 3804 2360 3832 2391
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4672 2400 4721 2428
rect 4672 2388 4678 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5868 2400 6377 2428
rect 5868 2388 5874 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7282 2388 7288 2440
rect 7340 2388 7346 2440
rect 7374 2388 7380 2440
rect 7432 2428 7438 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7432 2400 7665 2428
rect 7432 2388 7438 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 9140 2437 9168 2468
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 3292 2332 3832 2360
rect 3292 2320 3298 2332
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 3878 2292 3884 2304
rect 3467 2264 3884 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4580 2264 4905 2292
rect 4580 2252 4586 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7469 2295 7527 2301
rect 7469 2292 7481 2295
rect 6880 2264 7481 2292
rect 6880 2252 6886 2264
rect 7469 2261 7481 2264
rect 7515 2261 7527 2295
rect 7469 2255 7527 2261
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 7984 2264 8217 2292
rect 7984 2252 7990 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 1104 2202 10028 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 10028 2202
rect 1104 2128 10028 2150
<< via1 >>
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3884 10752 3936 10804
rect 4528 10752 4580 10804
rect 5264 10752 5316 10804
rect 5816 10752 5868 10804
rect 6460 10752 6512 10804
rect 7104 10752 7156 10804
rect 1952 10616 2004 10668
rect 2596 10616 2648 10668
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4620 10616 4672 10668
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8392 10616 8444 10668
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3240 10208 3292 10260
rect 4068 10208 4120 10260
rect 5264 10208 5316 10260
rect 2964 10072 3016 10124
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 4252 10115 4304 10124
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 5816 10208 5868 10260
rect 6184 10208 6236 10260
rect 6644 10208 6696 10260
rect 7564 10208 7616 10260
rect 7748 10208 7800 10260
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 2964 9979 3016 9988
rect 2964 9945 2973 9979
rect 2973 9945 3007 9979
rect 3007 9945 3016 9979
rect 2964 9936 3016 9945
rect 3516 10004 3568 10056
rect 4804 10004 4856 10056
rect 6184 10004 6236 10056
rect 3608 9936 3660 9988
rect 3332 9868 3384 9920
rect 4252 9868 4304 9920
rect 8208 10004 8260 10056
rect 6184 9868 6236 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2044 9664 2096 9716
rect 2964 9664 3016 9716
rect 3608 9664 3660 9716
rect 4436 9664 4488 9716
rect 4804 9664 4856 9716
rect 3516 9596 3568 9648
rect 3332 9528 3384 9580
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 5908 9120 5960 9172
rect 2688 9052 2740 9104
rect 5816 8984 5868 9036
rect 940 8848 992 8900
rect 5356 8916 5408 8968
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 4436 8848 4488 8900
rect 4620 8848 4672 8900
rect 3332 8780 3384 8832
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 3976 8780 4028 8832
rect 8024 8848 8076 8900
rect 4804 8780 4856 8832
rect 8668 8780 8720 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3424 8576 3476 8628
rect 3976 8508 4028 8560
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 4804 8440 4856 8492
rect 6276 8576 6328 8628
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 5172 8372 5224 8424
rect 5448 8440 5500 8492
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 7288 8576 7340 8628
rect 6828 8440 6880 8492
rect 5908 8372 5960 8424
rect 7288 8372 7340 8424
rect 7012 8304 7064 8356
rect 4712 8236 4764 8288
rect 5356 8236 5408 8288
rect 7104 8236 7156 8288
rect 7288 8236 7340 8288
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 7656 8279 7708 8288
rect 7656 8245 7665 8279
rect 7665 8245 7699 8279
rect 7699 8245 7708 8279
rect 7656 8236 7708 8245
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9220 8440 9272 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 9588 8347 9640 8356
rect 9588 8313 9597 8347
rect 9597 8313 9631 8347
rect 9631 8313 9640 8347
rect 9588 8304 9640 8313
rect 8668 8236 8720 8288
rect 9312 8236 9364 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 7012 8032 7064 8084
rect 4712 7964 4764 8016
rect 2320 7896 2372 7948
rect 3700 7896 3752 7948
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 4160 7828 4212 7880
rect 4620 7896 4672 7948
rect 5172 7896 5224 7948
rect 7380 7964 7432 8016
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 8208 8032 8260 8084
rect 9036 8032 9088 8084
rect 5448 7896 5500 7948
rect 6920 7896 6972 7948
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 5356 7828 5408 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 8116 7964 8168 8016
rect 3976 7760 4028 7812
rect 5448 7760 5500 7812
rect 5816 7760 5868 7812
rect 7104 7760 7156 7812
rect 8484 7828 8536 7880
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 9220 7828 9272 7880
rect 8208 7803 8260 7812
rect 8208 7769 8217 7803
rect 8217 7769 8251 7803
rect 8251 7769 8260 7803
rect 8208 7760 8260 7769
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4804 7692 4856 7744
rect 5172 7692 5224 7744
rect 8300 7692 8352 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 10140 7692 10192 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2136 7488 2188 7540
rect 3792 7488 3844 7540
rect 3976 7488 4028 7540
rect 3424 7420 3476 7472
rect 6644 7488 6696 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 7012 7488 7064 7540
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 8944 7488 8996 7540
rect 9128 7488 9180 7540
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 6552 7352 6604 7404
rect 6920 7420 6972 7472
rect 7472 7463 7524 7472
rect 7472 7429 7481 7463
rect 7481 7429 7515 7463
rect 7515 7429 7524 7463
rect 7472 7420 7524 7429
rect 5264 7284 5316 7336
rect 8116 7352 8168 7404
rect 8300 7352 8352 7404
rect 7840 7327 7892 7336
rect 6644 7216 6696 7268
rect 7196 7216 7248 7268
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 8024 7284 8076 7336
rect 4896 7148 4948 7200
rect 5356 7148 5408 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 7840 6944 7892 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8944 6987 8996 6996
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 4896 6876 4948 6928
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 4804 6808 4856 6860
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 3424 6740 3476 6792
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 3332 6715 3384 6724
rect 3332 6681 3341 6715
rect 3341 6681 3375 6715
rect 3375 6681 3384 6715
rect 3332 6672 3384 6681
rect 4068 6672 4120 6724
rect 4620 6740 4672 6792
rect 6460 6740 6512 6792
rect 7656 6740 7708 6792
rect 8576 6740 8628 6792
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 4712 6672 4764 6724
rect 3424 6647 3476 6656
rect 3424 6613 3439 6647
rect 3439 6613 3473 6647
rect 3473 6613 3476 6647
rect 3424 6604 3476 6613
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 6368 6647 6420 6656
rect 6368 6613 6377 6647
rect 6377 6613 6411 6647
rect 6411 6613 6420 6647
rect 6368 6604 6420 6613
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 3700 6400 3752 6452
rect 4620 6400 4672 6452
rect 5264 6400 5316 6452
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 6460 6400 6512 6452
rect 8484 6400 8536 6452
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 3976 6332 4028 6384
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 4804 6332 4856 6384
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 4620 6196 4672 6248
rect 5080 6196 5132 6248
rect 5540 6264 5592 6316
rect 6644 6264 6696 6316
rect 6920 6264 6972 6316
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 6460 6239 6512 6248
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 6920 6171 6972 6180
rect 6920 6137 6929 6171
rect 6929 6137 6963 6171
rect 6963 6137 6972 6171
rect 6920 6128 6972 6137
rect 7380 6128 7432 6180
rect 10140 6196 10192 6248
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 5448 6060 5500 6112
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 9036 6128 9088 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3608 5856 3660 5908
rect 4712 5856 4764 5908
rect 3056 5720 3108 5772
rect 2228 5652 2280 5704
rect 4804 5831 4856 5840
rect 4804 5797 4813 5831
rect 4813 5797 4847 5831
rect 4847 5797 4856 5831
rect 4804 5788 4856 5797
rect 6460 5856 6512 5908
rect 6644 5856 6696 5908
rect 8484 5856 8536 5908
rect 5816 5720 5868 5772
rect 4620 5652 4672 5704
rect 4804 5652 4856 5704
rect 5448 5695 5500 5704
rect 2872 5584 2924 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 5080 5627 5132 5636
rect 5080 5593 5089 5627
rect 5089 5593 5123 5627
rect 5123 5593 5132 5627
rect 5080 5584 5132 5593
rect 6184 5584 6236 5636
rect 8944 5788 8996 5840
rect 8300 5720 8352 5772
rect 9680 5720 9732 5772
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 9036 5652 9088 5704
rect 6276 5516 6328 5568
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 7196 5516 7248 5568
rect 9588 5584 9640 5636
rect 8024 5516 8076 5568
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2872 5312 2924 5364
rect 3056 5312 3108 5364
rect 3516 5312 3568 5364
rect 7380 5312 7432 5364
rect 8116 5312 8168 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 6368 5244 6420 5296
rect 6920 5244 6972 5296
rect 7196 5244 7248 5296
rect 7656 5287 7708 5296
rect 7656 5253 7665 5287
rect 7665 5253 7699 5287
rect 7699 5253 7708 5287
rect 7656 5244 7708 5253
rect 3332 5176 3384 5228
rect 4068 5176 4120 5228
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 5264 5108 5316 5160
rect 5632 5040 5684 5092
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 6276 5176 6328 5228
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 8484 5244 8536 5296
rect 8852 5244 8904 5296
rect 8300 5108 8352 5160
rect 4988 4972 5040 5024
rect 5264 4972 5316 5024
rect 6092 4972 6144 5024
rect 8208 4972 8260 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2136 4768 2188 4820
rect 3056 4768 3108 4820
rect 4896 4768 4948 4820
rect 5448 4768 5500 4820
rect 6092 4768 6144 4820
rect 3424 4700 3476 4752
rect 6276 4700 6328 4752
rect 4988 4632 5040 4684
rect 8300 4632 8352 4684
rect 8760 4632 8812 4684
rect 9496 4632 9548 4684
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 4620 4564 4672 4616
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 2136 4496 2188 4548
rect 3976 4428 4028 4480
rect 4804 4428 4856 4480
rect 8668 4428 8720 4480
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9496 4471 9548 4480
rect 9496 4437 9505 4471
rect 9505 4437 9539 4471
rect 9539 4437 9548 4471
rect 9496 4428 9548 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2136 4267 2188 4276
rect 2136 4233 2145 4267
rect 2145 4233 2179 4267
rect 2179 4233 2188 4267
rect 2136 4224 2188 4233
rect 4804 4224 4856 4276
rect 5264 4224 5316 4276
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 3056 4088 3108 4140
rect 3424 4088 3476 4140
rect 6460 4088 6512 4140
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 5540 4020 5592 4072
rect 9496 4088 9548 4140
rect 2412 3927 2464 3936
rect 2412 3893 2421 3927
rect 2421 3893 2455 3927
rect 2455 3893 2464 3927
rect 2412 3884 2464 3893
rect 9588 3927 9640 3936
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3608 3680 3660 3732
rect 4620 3680 4672 3732
rect 3056 3544 3108 3596
rect 4712 3544 4764 3596
rect 5540 3476 5592 3528
rect 1584 3408 1636 3460
rect 2412 3408 2464 3460
rect 7564 3451 7616 3460
rect 7564 3417 7573 3451
rect 7573 3417 7607 3451
rect 7607 3417 7616 3451
rect 7564 3408 7616 3417
rect 7472 3340 7524 3392
rect 7840 3383 7892 3392
rect 7840 3349 7849 3383
rect 7849 3349 7883 3383
rect 7883 3349 7892 3383
rect 7840 3340 7892 3349
rect 7932 3340 7984 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 7564 3179 7616 3188
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 6644 3068 6696 3120
rect 7564 3145 7573 3179
rect 7573 3145 7607 3179
rect 7607 3145 7616 3179
rect 7564 3136 7616 3145
rect 7840 3136 7892 3188
rect 7196 3068 7248 3120
rect 7932 3068 7984 3120
rect 4160 2932 4212 2984
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 7472 3000 7524 3052
rect 7564 3000 7616 3052
rect 4988 2864 5040 2916
rect 7104 2932 7156 2984
rect 7196 2907 7248 2916
rect 3700 2796 3752 2848
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 6000 2796 6052 2848
rect 7196 2873 7205 2907
rect 7205 2873 7239 2907
rect 7239 2873 7248 2907
rect 7196 2864 7248 2873
rect 7380 2796 7432 2848
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 9680 2796 9732 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 4804 2592 4856 2644
rect 6644 2592 6696 2644
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 6000 2456 6052 2508
rect 7104 2524 7156 2576
rect 3700 2388 3752 2440
rect 3240 2320 3292 2372
rect 4620 2388 4672 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5816 2388 5868 2440
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7380 2388 7432 2440
rect 7748 2388 7800 2440
rect 8392 2388 8444 2440
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 3884 2252 3936 2304
rect 4528 2252 4580 2304
rect 6828 2252 6880 2304
rect 7932 2252 7984 2304
rect 8392 2252 8444 2304
rect 9036 2252 9088 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 1950 12517 2006 13317
rect 2594 12517 2650 13317
rect 3238 12517 3294 13317
rect 3882 12517 3938 13317
rect 4526 12517 4582 13317
rect 5170 12517 5226 13317
rect 5814 12517 5870 13317
rect 6458 12517 6514 13317
rect 7102 12517 7158 13317
rect 7746 12517 7802 13317
rect 8390 12517 8446 13317
rect 1964 10674 1992 12517
rect 2608 10674 2636 12517
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2056 9722 2084 10542
rect 2976 10130 3004 10542
rect 3252 10266 3280 12517
rect 3896 10810 3924 12517
rect 4540 10810 4568 12517
rect 5184 11098 5212 12517
rect 5184 11070 5304 11098
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10810 5304 11070
rect 5828 10810 5856 12517
rect 6472 10810 6500 12517
rect 7116 10810 7144 12517
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 4080 10266 4108 10610
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4632 10130 4660 10610
rect 5276 10266 5304 10610
rect 5828 10266 5856 10610
rect 6656 10266 6684 10610
rect 7576 10266 7604 10610
rect 7760 10266 7788 12517
rect 8404 10674 8432 12517
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9722 3004 9930
rect 3344 9926 3372 10066
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3344 9586 3372 9862
rect 3528 9654 3556 9998
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3620 9722 3648 9930
rect 4264 9926 4292 10066
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4448 9722 4476 10066
rect 6196 10062 6224 10202
rect 8220 10062 8248 10542
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 4816 9722 4844 9998
rect 6196 9926 6224 9998
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3620 9518 3648 9658
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 938 8936 994 8945
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 940 8842 992 8848
rect 2700 8498 2728 9046
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 7954 2360 8366
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7546 2176 7822
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 3344 7410 3372 8774
rect 3436 8634 3464 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3436 7478 3464 8570
rect 3988 8566 4016 8774
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3344 6730 3372 7346
rect 3436 6798 3464 7414
rect 3712 7410 3740 7890
rect 3988 7818 4016 8502
rect 4448 8412 4476 8842
rect 4632 8514 4660 8842
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4632 8486 4752 8514
rect 4816 8498 4844 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4448 8384 4660 8412
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8384
rect 4724 8294 4752 8486
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 8022 4752 8230
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4618 7848 4674 7857
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7546 3832 7686
rect 3988 7546 4016 7754
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3424 6792 3476 6798
rect 3608 6792 3660 6798
rect 3476 6740 3556 6746
rect 3424 6734 3556 6740
rect 3608 6734 3660 6740
rect 3332 6724 3384 6730
rect 3436 6718 3556 6734
rect 3332 6666 3384 6672
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6322 3464 6598
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5710 2268 6054
rect 3068 5778 3096 6258
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1398 4176 1454 4185
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 1400 4082 1452 4088
rect 1596 3466 1624 5510
rect 2884 5370 2912 5578
rect 3068 5370 3096 5714
rect 3528 5370 3556 6718
rect 3620 5914 3648 6734
rect 3712 6458 3740 7346
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3988 6390 4016 7482
rect 4172 7290 4200 7822
rect 4618 7783 4674 7792
rect 4080 7262 4200 7290
rect 4080 6882 4108 7262
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4080 6866 4384 6882
rect 4080 6860 4396 6866
rect 4080 6854 4344 6860
rect 4344 6802 4396 6808
rect 4632 6798 4660 7783
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4724 6730 4752 7958
rect 4816 7750 4844 8434
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5184 7954 5212 8366
rect 5368 8294 5396 8910
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5460 7954 5488 8434
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5184 7750 5212 7890
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 4816 6866 4844 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6934 4936 7142
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2148 4826 2176 5102
rect 3068 4826 3096 5306
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 2148 4282 2176 4490
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 3068 4146 3096 4762
rect 3344 4622 3372 5170
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3436 4146 3464 4694
rect 3528 4622 3556 5306
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3466 2452 3878
rect 3068 3602 3096 4082
rect 3620 3738 3648 4558
rect 3988 4486 4016 6326
rect 4080 5234 4108 6666
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6458 4660 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6458 5304 7278
rect 5368 7206 5396 7822
rect 5828 7818 5856 8978
rect 5920 8430 5948 9114
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 6288 8634 6316 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 4804 6384 4856 6390
rect 5460 6338 5488 7754
rect 6472 6798 6500 8434
rect 6840 7546 6868 8434
rect 6932 7954 6960 8910
rect 7300 8634 7328 8910
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7470 8392 7526 8401
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7024 8090 7052 8298
rect 7300 8294 7328 8366
rect 7470 8327 7526 8336
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7024 7546 7052 8026
rect 7116 7818 7144 8230
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 4804 6326 4856 6332
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5710 4660 6190
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3738 4660 4558
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4724 3602 4752 5850
rect 4816 5846 4844 6326
rect 5368 6322 5580 6338
rect 5356 6316 5592 6322
rect 5408 6310 5540 6316
rect 5356 6258 5408 6264
rect 5540 6258 5592 6264
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4816 5710 4844 5782
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 4842 4844 5646
rect 5092 5642 5120 6190
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5368 5234 5396 6258
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 5710 5488 6054
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5264 5160 5316 5166
rect 5316 5108 5396 5114
rect 5264 5102 5396 5108
rect 5276 5086 5396 5102
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 4816 4826 4936 4842
rect 4816 4820 4948 4826
rect 4816 4814 4896 4820
rect 4896 4762 4948 4768
rect 5000 4690 5028 4966
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4282 4844 4422
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5276 4282 5304 4966
rect 5368 4282 5396 5086
rect 5460 4826 5488 5170
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5552 4078 5580 5170
rect 5644 5098 5672 6394
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6196 5234 6224 5578
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5234 6316 5510
rect 6380 5302 6408 6598
rect 6472 6458 6500 6734
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6564 6338 6592 7346
rect 6656 7274 6684 7482
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6472 6310 6592 6338
rect 6656 6322 6684 7210
rect 6932 6322 6960 7414
rect 7208 7274 7236 7890
rect 7300 7546 7328 8230
rect 7392 8022 7420 8230
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7484 7886 7512 8327
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 8022 7696 8230
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7484 7478 7512 7822
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 8036 7342 8064 8842
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8482 8392 8538 8401
rect 8482 8327 8538 8336
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7410 8156 7958
rect 8220 7818 8248 8026
rect 8496 7886 8524 8327
rect 8680 8294 8708 8774
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 9048 8090 9076 8434
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9232 7886 9260 8434
rect 9324 8401 9352 8434
rect 9310 8392 9366 8401
rect 9310 8327 9366 8336
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9312 8288 9364 8294
rect 9600 8265 9628 8298
rect 9312 8230 9364 8236
rect 9586 8256 9642 8265
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7410 8340 7686
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7852 7002 7880 7278
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 6644 6316 6696 6322
rect 6472 6254 6500 6310
rect 6644 6258 6696 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 5914 6500 6190
rect 6656 5914 6684 6258
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4826 6132 4966
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6288 4758 6316 5170
rect 6472 5166 6500 5510
rect 6932 5302 6960 6122
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5302 7236 5510
rect 7392 5370 7420 6122
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7668 5302 7696 6734
rect 8036 5574 8064 7278
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8312 5778 8340 6938
rect 8496 6458 8524 7822
rect 8588 6798 8616 7822
rect 9140 7546 9168 7822
rect 9324 7750 9352 8230
rect 9586 8191 9642 8200
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8956 7002 8984 7482
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9140 6798 9168 7482
rect 9324 6866 9352 7686
rect 10152 7585 10180 7686
rect 10138 7576 10194 7585
rect 10138 7511 10194 7520
rect 9586 6896 9642 6905
rect 9312 6860 9364 6866
rect 9586 6831 9642 6840
rect 9312 6802 9364 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 6458 9444 6734
rect 9600 6662 9628 6831
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8496 5914 8524 6190
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8128 5370 8156 5646
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 8312 5166 8340 5714
rect 8496 5302 8524 5850
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6472 4146 6500 5102
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4622 8248 4966
rect 8312 4690 8340 5102
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8680 4486 8708 6258
rect 8944 6248 8996 6254
rect 10140 6248 10192 6254
rect 8944 6190 8996 6196
rect 10138 6216 10140 6225
rect 10192 6216 10194 6225
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 4690 8800 5510
rect 8864 5302 8892 6054
rect 8956 5846 8984 6190
rect 9036 6180 9088 6186
rect 10138 6151 10194 6160
rect 9036 6122 9088 6128
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9048 5710 9076 6122
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9496 5568 9548 5574
rect 9600 5545 9628 5578
rect 9496 5510 9548 5516
rect 9586 5536 9642 5545
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 9508 4690 9536 5510
rect 9586 5471 9642 5480
rect 9692 5370 9720 5714
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9586 4856 9642 4865
rect 9586 4791 9642 4800
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 9232 4282 9260 4558
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 8850 4176 8906 4185
rect 6460 4140 6512 4146
rect 9508 4146 9536 4422
rect 8850 4111 8852 4120
rect 6460 4082 6512 4088
rect 8904 4111 8906 4120
rect 9496 4140 9548 4146
rect 8852 4082 8904 4088
rect 9496 4082 9548 4088
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 5552 3534 5580 4014
rect 9600 3942 9628 4791
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 1584 3460 1636 3466
rect 1584 3402 1636 3408
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 4160 2984 4212 2990
rect 4080 2932 4160 2938
rect 4080 2926 4212 2932
rect 4080 2910 4200 2926
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2446 3740 2790
rect 4080 2514 4108 2910
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4632 2446 4660 2790
rect 4816 2650 4844 2994
rect 5000 2922 5028 2994
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 6012 2854 6040 2994
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 6012 2514 6040 2790
rect 6656 2650 6684 3062
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7116 2774 7144 2926
rect 7208 2922 7236 3062
rect 7484 3058 7512 3334
rect 7576 3194 7604 3402
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7852 3194 7880 3334
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7576 3058 7604 3130
rect 7944 3126 7972 3334
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 7116 2746 7328 2774
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3252 800 3280 2314
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 3896 800 3924 2246
rect 4540 800 4568 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2382
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 5828 800 5856 2382
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6472 870 6592 898
rect 6472 800 6500 870
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 6564 762 6592 870
rect 6840 762 6868 2246
rect 7116 800 7144 2518
rect 7300 2446 7328 2746
rect 7392 2446 7420 2790
rect 7760 2446 7788 2790
rect 8404 2446 8432 2790
rect 8496 2446 8524 2790
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 7932 2304 7984 2310
rect 7760 2264 7932 2292
rect 7760 800 7788 2264
rect 7932 2246 7984 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 8404 800 8432 2246
rect 9048 800 9076 2246
rect 9692 800 9720 2790
rect 6564 734 6868 762
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
<< via2 >>
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 4618 7792 4674 7848
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 7470 8336 7526 8392
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 8482 8336 8538 8392
rect 9310 8336 9366 8392
rect 9586 8200 9642 8256
rect 10138 7520 10194 7576
rect 9586 6840 9642 6896
rect 10138 6196 10140 6216
rect 10140 6196 10192 6216
rect 10192 6196 10194 6216
rect 10138 6160 10194 6196
rect 9586 5480 9642 5536
rect 9586 4800 9642 4856
rect 8850 4140 8906 4176
rect 8850 4120 8852 4140
rect 8852 4120 8904 4140
rect 8904 4120 8906 4140
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 7465 8394 7531 8397
rect 8477 8394 8543 8397
rect 9305 8394 9371 8397
rect 7465 8392 9371 8394
rect 7465 8336 7470 8392
rect 7526 8336 8482 8392
rect 8538 8336 9310 8392
rect 9366 8336 9371 8392
rect 7465 8334 9371 8336
rect 7465 8331 7531 8334
rect 8477 8331 8543 8334
rect 9305 8331 9371 8334
rect 0 8258 800 8288
rect 9581 8258 9647 8261
rect 10373 8258 11173 8288
rect 0 8198 2330 8258
rect 0 8168 800 8198
rect 2270 7850 2330 8198
rect 9581 8256 11173 8258
rect 9581 8200 9586 8256
rect 9642 8200 11173 8256
rect 9581 8198 11173 8200
rect 9581 8195 9647 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 10373 8168 11173 8198
rect 4210 8127 4526 8128
rect 4613 7850 4679 7853
rect 2270 7848 4679 7850
rect 2270 7792 4618 7848
rect 4674 7792 4679 7848
rect 2270 7790 4679 7792
rect 4613 7787 4679 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 10133 7578 10199 7581
rect 10373 7578 11173 7608
rect 10133 7576 11173 7578
rect 10133 7520 10138 7576
rect 10194 7520 11173 7576
rect 10133 7518 11173 7520
rect 10133 7515 10199 7518
rect 10373 7488 11173 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 9581 6898 9647 6901
rect 10373 6898 11173 6928
rect 9581 6896 11173 6898
rect 9581 6840 9586 6896
rect 9642 6840 11173 6896
rect 9581 6838 11173 6840
rect 9581 6835 9647 6838
rect 10373 6808 11173 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 10133 6218 10199 6221
rect 10373 6218 11173 6248
rect 10133 6216 11173 6218
rect 10133 6160 10138 6216
rect 10194 6160 11173 6216
rect 10133 6158 11173 6160
rect 10133 6155 10199 6158
rect 10373 6128 11173 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 9581 5538 9647 5541
rect 10373 5538 11173 5568
rect 9581 5536 11173 5538
rect 9581 5480 9586 5536
rect 9642 5480 11173 5536
rect 9581 5478 11173 5480
rect 9581 5475 9647 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 10373 5448 11173 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 9581 4858 9647 4861
rect 10373 4858 11173 4888
rect 9581 4856 11173 4858
rect 9581 4800 9586 4856
rect 9642 4800 11173 4856
rect 9581 4798 11173 4800
rect 9581 4795 9647 4798
rect 10373 4768 11173 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 8845 4178 8911 4181
rect 10373 4178 11173 4208
rect 8845 4176 11173 4178
rect 8845 4120 8850 4176
rect 8906 4120 11173 4176
rect 8845 4118 11173 4120
rect 8845 4115 8911 4118
rect 10373 4088 11173 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 10368 4528 10928
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 10928
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _043_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _044_
timestamp 1707688321
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _045_
timestamp 1707688321
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _046_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _047_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 5336 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 4784 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _049_
timestamp 1707688321
transform 1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _050_
timestamp 1707688321
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _051_
timestamp 1707688321
transform 1 0 4784 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _052_
timestamp 1707688321
transform -1 0 9384 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 8924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4600 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _057_
timestamp 1707688321
transform 1 0 4048 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 7820 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _059_
timestamp 1707688321
transform -1 0 6256 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _060_
timestamp 1707688321
transform 1 0 7176 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _061_
timestamp 1707688321
transform 1 0 6532 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8924 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _063_
timestamp 1707688321
transform -1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _064_
timestamp 1707688321
transform -1 0 3680 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _065_
timestamp 1707688321
transform 1 0 3404 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _066_
timestamp 1707688321
transform 1 0 6348 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _067_
timestamp 1707688321
transform -1 0 4692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _068_
timestamp 1707688321
transform 1 0 5704 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _069_
timestamp 1707688321
transform 1 0 5060 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _070_
timestamp 1707688321
transform 1 0 6992 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _073_
timestamp 1707688321
transform 1 0 8464 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6992 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _077_
timestamp 1707688321
transform -1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _078_
timestamp 1707688321
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4324 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _080_
timestamp 1707688321
transform -1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _081_
timestamp 1707688321
transform -1 0 4692 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 5428 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _083_
timestamp 1707688321
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _085_
timestamp 1707688321
transform -1 0 4324 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _086_
timestamp 1707688321
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 4600 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _088_
timestamp 1707688321
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _089_
timestamp 1707688321
transform 1 0 5152 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _090_
timestamp 1707688321
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _091_
timestamp 1707688321
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _092_
timestamp 1707688321
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _093_
timestamp 1707688321
transform -1 0 7728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _094_
timestamp 1707688321
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _095_
timestamp 1707688321
transform -1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 6900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _097_
timestamp 1707688321
transform 1 0 8188 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 8832 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _099_
timestamp 1707688321
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _100_
timestamp 1707688321
transform 1 0 6440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 7912 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _102_
timestamp 1707688321
transform 1 0 6808 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 7268 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1707688321
transform -1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1748 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _107_
timestamp 1707688321
transform 1 0 2300 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _108_
timestamp 1707688321
transform -1 0 6716 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _109_
timestamp 1707688321
transform 1 0 3680 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _110_
timestamp 1707688321
transform 1 0 3036 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _111_
timestamp 1707688321
transform 1 0 3128 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _112_
timestamp 1707688321
transform 1 0 4692 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _113_
timestamp 1707688321
transform -1 0 8648 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _114_
timestamp 1707688321
transform -1 0 8556 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _115_
timestamp 1707688321
transform 1 0 6900 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _116_
timestamp 1707688321
transform 1 0 7820 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _117_
timestamp 1707688321
transform -1 0 7268 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _118_
timestamp 1707688321
transform 1 0 1748 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _118__34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _119__35
timestamp 1707688321
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1380 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 1707688321
transform -1 0 3220 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 1707688321
transform 1 0 7912 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_osc_ck $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5060 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_osc_ck
timestamp 1707688321
transform -1 0 4692 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_osc_ck
timestamp 1707688321
transform 1 0 6992 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1707688321
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_79
timestamp 1707688321
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1707688321
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1707688321
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1707688321
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_31
timestamp 1707688321
transform 1 0 3956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5152 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1707688321
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_85
timestamp 1707688321
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_89
timestamp 1707688321
transform 1 0 9292 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_23
timestamp 1707688321
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1707688321
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1707688321
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_38
timestamp 1707688321
transform 1 0 4600 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_50
timestamp 1707688321
transform 1 0 5704 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_62
timestamp 1707688321
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_74
timestamp 1707688321
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1707688321
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1707688321
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_93
timestamp 1707688321
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_6
timestamp 1707688321
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_16
timestamp 1707688321
transform 1 0 2576 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_43
timestamp 1707688321
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_48
timestamp 1707688321
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1707688321
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1707688321
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_81
timestamp 1707688321
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_23
timestamp 1707688321
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_37
timestamp 1707688321
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_60
timestamp 1707688321
transform 1 0 6624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1707688321
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_92
timestamp 1707688321
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1707688321
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_39
timestamp 1707688321
transform 1 0 4692 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_72
timestamp 1707688321
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_6
timestamp 1707688321
transform 1 0 1656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1707688321
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_55
timestamp 1707688321
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_92
timestamp 1707688321
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1707688321
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_11
timestamp 1707688321
transform 1 0 2116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_15
timestamp 1707688321
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1707688321
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_69
timestamp 1707688321
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_77
timestamp 1707688321
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1707688321
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_15
timestamp 1707688321
transform 1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_23
timestamp 1707688321
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_29
timestamp 1707688321
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_39
timestamp 1707688321
transform 1 0 4692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_63
timestamp 1707688321
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1707688321
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 1707688321
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_19
timestamp 1707688321
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 1707688321
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1707688321
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_71
timestamp 1707688321
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1707688321
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_37
timestamp 1707688321
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1707688321
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_11
timestamp 1707688321
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 1707688321
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1707688321
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1707688321
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_75
timestamp 1707688321
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_7
timestamp 1707688321
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_19
timestamp 1707688321
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1707688321
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_61
timestamp 1707688321
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1707688321
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_93
timestamp 1707688321
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1707688321
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_15
timestamp 1707688321
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_23
timestamp 1707688321
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_31
timestamp 1707688321
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 1707688321
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1707688321
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1707688321
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1707688321
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1707688321
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_93
timestamp 1707688321
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1707688321
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_15
timestamp 1707688321
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1707688321
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_69
timestamp 1707688321
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 1707688321
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1707688321
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1707688321
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1707688321
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1707688321
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_27
timestamp 1707688321
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_29
timestamp 1707688321
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_37
timestamp 1707688321
transform 1 0 4508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1707688321
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1707688321
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_72
timestamp 1707688321
transform 1 0 7728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_85
timestamp 1707688321
transform 1 0 8924 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_93
timestamp 1707688321
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1707688321
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1707688321
transform 1 0 5428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1707688321
transform -1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1707688321
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1707688321
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1707688321
transform -1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1707688321
transform 1 0 5244 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1707688321
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1707688321
transform 1 0 7912 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1707688321
transform 1 0 1748 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1707688321
transform 1 0 2668 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1707688321
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1707688321
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1707688321
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1707688321
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1707688321
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1707688321
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1707688321
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1707688321
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1707688321
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1707688321
transform 1 0 9384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1707688321
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1707688321
transform 1 0 5152 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1707688321
transform 1 0 3956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1707688321
transform -1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1707688321
transform 1 0 7820 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1707688321
transform 1 0 4600 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1707688321
transform 1 0 6532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1707688321
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1707688321
transform -1 0 7728 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_16
timestamp 1707688321
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1707688321
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_17
timestamp 1707688321
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1707688321
transform -1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_18
timestamp 1707688321
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1707688321
transform -1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_19
timestamp 1707688321
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1707688321
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_20
timestamp 1707688321
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1707688321
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_21
timestamp 1707688321
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1707688321
transform -1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_22
timestamp 1707688321
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1707688321
transform -1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_23
timestamp 1707688321
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1707688321
transform -1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_24
timestamp 1707688321
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1707688321
transform -1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_25
timestamp 1707688321
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1707688321
transform -1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_26
timestamp 1707688321
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1707688321
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_27
timestamp 1707688321
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1707688321
transform -1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_28
timestamp 1707688321
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1707688321
transform -1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_29
timestamp 1707688321
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1707688321
transform -1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_30
timestamp 1707688321
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1707688321
transform -1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_31
timestamp 1707688321
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1707688321
transform -1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp 1707688321
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 1707688321
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_35
timestamp 1707688321
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 1707688321
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 1707688321
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_38
timestamp 1707688321
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_39
timestamp 1707688321
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_40
timestamp 1707688321
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_41
timestamp 1707688321
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_42
timestamp 1707688321
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_43
timestamp 1707688321
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_44
timestamp 1707688321
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_45
timestamp 1707688321
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_46
timestamp 1707688321
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_47
timestamp 1707688321
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_48
timestamp 1707688321
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_49
timestamp 1707688321
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_50
timestamp 1707688321
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_51
timestamp 1707688321
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_52
timestamp 1707688321
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_53
timestamp 1707688321
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_54
timestamp 1707688321
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_55
timestamp 1707688321
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_56
timestamp 1707688321
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_57
timestamp 1707688321
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1707688321
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 10928 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 10928 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 brout_filt
port 3 nsew signal input
flabel metal3 s 10373 6128 11173 6248 0 FreeSans 480 0 0 0 dcomp
port 4 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 ena
port 5 nsew signal input
flabel metal3 s 10373 4088 11173 4208 0 FreeSans 480 0 0 0 force_dis_rc_osc
port 6 nsew signal input
flabel metal3 s 10373 5448 11173 5568 0 FreeSans 480 0 0 0 force_ena_rc_osc
port 7 nsew signal input
flabel metal3 s 10373 7488 11173 7608 0 FreeSans 480 0 0 0 force_short_oneshot
port 8 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 osc_ck
port 9 nsew signal input
flabel metal3 s 10373 4768 11173 4888 0 FreeSans 480 0 0 0 osc_ena
port 16 nsew signal output
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 otrip[0]
port 10 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 otrip[1]
port 11 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 otrip[2]
port 12 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 otrip_decoded[0]
port 17 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 otrip_decoded[1]
port 18 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 otrip_decoded[2]
port 19 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 otrip_decoded[3]
port 20 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 otrip_decoded[4]
port 21 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 otrip_decoded[5]
port 22 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 otrip_decoded[6]
port 23 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 otrip_decoded[7]
port 24 nsew signal output
flabel metal3 s 10373 6808 11173 6928 0 FreeSans 480 0 0 0 outb_unbuf
port 25 nsew signal output
flabel metal3 s 10373 8168 11173 8288 0 FreeSans 480 0 0 0 timed_out
port 26 nsew signal output
flabel metal2 s 8390 12517 8446 13317 0 FreeSans 224 90 0 0 vtrip[0]
port 13 nsew signal input
flabel metal2 s 1950 12517 2006 13317 0 FreeSans 224 90 0 0 vtrip[1]
port 14 nsew signal input
flabel metal2 s 2594 12517 2650 13317 0 FreeSans 224 90 0 0 vtrip[2]
port 15 nsew signal input
flabel metal2 s 5170 12517 5226 13317 0 FreeSans 224 90 0 0 vtrip_decoded[0]
port 27 nsew signal output
flabel metal2 s 3882 12517 3938 13317 0 FreeSans 224 90 0 0 vtrip_decoded[1]
port 28 nsew signal output
flabel metal2 s 3238 12517 3294 13317 0 FreeSans 224 90 0 0 vtrip_decoded[2]
port 29 nsew signal output
flabel metal2 s 7746 12517 7802 13317 0 FreeSans 224 90 0 0 vtrip_decoded[3]
port 30 nsew signal output
flabel metal2 s 4526 12517 4582 13317 0 FreeSans 224 90 0 0 vtrip_decoded[4]
port 31 nsew signal output
flabel metal2 s 6458 12517 6514 13317 0 FreeSans 224 90 0 0 vtrip_decoded[5]
port 32 nsew signal output
flabel metal2 s 5814 12517 5870 13317 0 FreeSans 224 90 0 0 vtrip_decoded[6]
port 33 nsew signal output
flabel metal2 s 7102 12517 7158 13317 0 FreeSans 224 90 0 0 vtrip_decoded[7]
port 34 nsew signal output
rlabel metal1 5566 10880 5566 10880 0 VGND
rlabel metal1 5566 10336 5566 10336 0 VPWR
rlabel metal2 2438 3672 2438 3672 0 _000_
rlabel metal2 2162 4386 2162 4386 0 _001_
rlabel metal2 2162 7684 2162 7684 0 _002_
rlabel metal2 2714 8772 2714 8772 0 _003_
rlabel metal1 5746 8602 5746 8602 0 _004_
rlabel metal1 3910 7310 3910 7310 0 _005_
rlabel metal2 3450 6460 3450 6460 0 _006_
rlabel metal1 3496 4114 3496 4114 0 _007_
rlabel metal1 5060 4658 5060 4658 0 _008_
rlabel metal2 8234 4794 8234 4794 0 _009_
rlabel metal1 7544 5066 7544 5066 0 _010_
rlabel metal1 8096 8602 8096 8602 0 _011_
rlabel metal1 8280 7378 8280 7378 0 _012_
rlabel metal1 7084 7854 7084 7854 0 _013_
rlabel metal1 5152 6426 5152 6426 0 _014_
rlabel metal1 4278 5712 4278 5712 0 _015_
rlabel metal1 3772 5882 3772 5882 0 _016_
rlabel metal1 3864 3706 3864 3706 0 _017_
rlabel metal1 5290 4182 5290 4182 0 _018_
rlabel metal2 5382 4675 5382 4675 0 _019_
rlabel metal1 7176 5134 7176 5134 0 _020_
rlabel metal1 6992 5202 6992 5202 0 _021_
rlabel metal1 8878 8398 8878 8398 0 _022_
rlabel metal1 9016 8330 9016 8330 0 _023_
rlabel metal1 8142 7888 8142 7888 0 _024_
rlabel metal1 7958 7820 7958 7820 0 _025_
rlabel metal1 7498 7990 7498 7990 0 _026_
rlabel metal2 7682 8126 7682 8126 0 _027_
rlabel metal1 8878 8058 8878 8058 0 _028_
rlabel metal2 9246 4420 9246 4420 0 _029_
rlabel metal1 5060 8330 5060 8330 0 _030_
rlabel via1 5382 6307 5382 6307 0 _031_
rlabel metal1 4646 5882 4646 5882 0 _032_
rlabel metal1 6394 5644 6394 5644 0 _033_
rlabel metal2 6486 4624 6486 4624 0 _034_
rlabel metal2 6486 6052 6486 6052 0 _035_
rlabel metal1 8142 7514 8142 7514 0 _036_
rlabel metal1 9430 4658 9430 4658 0 _037_
rlabel metal1 3496 7446 3496 7446 0 _038_
rlabel viali 5838 8466 5838 8466 0 _039_
rlabel metal1 5566 8262 5566 8262 0 _040_
rlabel metal1 4968 8398 4968 8398 0 _041_
rlabel metal1 4937 6290 4937 6290 0 _042_
rlabel metal3 1050 4148 1050 4148 0 brout_filt
rlabel metal2 6394 5950 6394 5950 0 clknet_0_osc_ck
rlabel metal2 2346 8160 2346 8160 0 clknet_1_0__leaf_osc_ck
rlabel metal1 6808 8942 6808 8942 0 clknet_1_1__leaf_osc_ck
rlabel metal1 5198 5678 5198 5678 0 clr_cnt
rlabel metal1 1794 4794 1794 4794 0 clr_cnt_sb
rlabel metal1 3910 3638 3910 3638 0 clr_cnt_sb_stg1
rlabel metal1 5152 7718 5152 7718 0 cnt\[0\]
rlabel metal1 9407 7514 9407 7514 0 cnt\[10\]
rlabel metal1 6946 8330 6946 8330 0 cnt\[11\]
rlabel metal1 4439 8262 4439 8262 0 cnt\[1\]
rlabel metal1 4876 7718 4876 7718 0 cnt\[2\]
rlabel metal1 5221 7174 5221 7174 0 cnt\[3\]
rlabel metal1 5451 6358 5451 6358 0 cnt\[4\]
rlabel metal2 5566 4352 5566 4352 0 cnt\[5\]
rlabel metal1 6072 5202 6072 5202 0 cnt\[6\]
rlabel metal1 6440 5202 6440 5202 0 cnt\[7\]
rlabel metal1 6624 6290 6624 6290 0 cnt\[8\]
rlabel metal2 9338 7276 9338 7276 0 cnt\[9\]
rlabel metal1 9706 6256 9706 6256 0 dcomp
rlabel metal2 8878 5678 8878 5678 0 dcomp_ena_rsb
rlabel metal1 9108 5746 9108 5746 0 dcomp_retimed
rlabel metal3 820 8908 820 8908 0 ena
rlabel via2 8878 4131 8878 4131 0 force_dis_rc_osc
rlabel metal1 8602 5644 8602 5644 0 force_ena_rc_osc
rlabel metal1 9936 7854 9936 7854 0 force_short_oneshot
rlabel metal1 1932 4114 1932 4114 0 net1
rlabel metal1 7741 9894 7741 9894 0 net10
rlabel metal1 3818 9588 3818 9588 0 net11
rlabel metal1 3542 9554 3542 9554 0 net12
rlabel metal1 9476 4114 9476 4114 0 net13
rlabel metal1 9430 3094 9430 3094 0 net14
rlabel metal1 4692 2414 4692 2414 0 net15
rlabel metal1 3680 2414 3680 2414 0 net16
rlabel metal1 9154 2448 9154 2448 0 net17
rlabel metal2 7314 2587 7314 2587 0 net18
rlabel metal1 7912 2414 7912 2414 0 net19
rlabel metal2 8510 5746 8510 5746 0 net2
rlabel metal1 7544 2414 7544 2414 0 net20
rlabel metal2 8510 2618 8510 2618 0 net21
rlabel metal2 9430 6596 9430 6596 0 net22
rlabel metal1 9384 8466 9384 8466 0 net23
rlabel metal1 5152 10234 5152 10234 0 net24
rlabel metal1 3864 10234 3864 10234 0 net25
rlabel metal1 3220 9690 3220 9690 0 net26
rlabel metal1 7728 9962 7728 9962 0 net27
rlabel metal2 4646 10370 4646 10370 0 net28
rlabel metal1 6486 10234 6486 10234 0 net29
rlabel metal1 3818 8874 3818 8874 0 net3
rlabel metal1 5750 10234 5750 10234 0 net30
rlabel metal1 7498 10234 7498 10234 0 net31
rlabel metal2 6486 7616 6486 7616 0 net32
rlabel metal1 7919 4522 7919 4522 0 net33
rlabel metal1 2208 5678 2208 5678 0 net34
rlabel metal1 1656 3434 1656 3434 0 net35
rlabel metal2 2898 5474 2898 5474 0 net36
rlabel metal1 2898 4488 2898 4488 0 net37
rlabel metal1 7268 5270 7268 5270 0 net38
rlabel metal1 3496 7514 3496 7514 0 net39
rlabel metal1 9108 4114 9108 4114 0 net4
rlabel metal1 8924 4658 8924 4658 0 net5
rlabel metal1 6670 7412 6670 7412 0 net6
rlabel metal1 4232 2958 4232 2958 0 net7
rlabel metal1 4646 3026 4646 3026 0 net8
rlabel metal1 4646 2958 4646 2958 0 net9
rlabel metal3 1487 8228 1487 8228 0 osc_ck
rlabel metal2 9614 4369 9614 4369 0 osc_ena
rlabel metal2 3266 1554 3266 1554 0 otrip[0]
rlabel metal2 5198 1027 5198 1027 0 otrip[1]
rlabel metal2 5842 1588 5842 1588 0 otrip[2]
rlabel metal1 9660 2822 9660 2822 0 otrip_decoded[0]
rlabel metal2 4554 1520 4554 1520 0 otrip_decoded[1]
rlabel metal2 3910 1520 3910 1520 0 otrip_decoded[2]
rlabel metal2 9062 1520 9062 1520 0 otrip_decoded[3]
rlabel metal2 6486 823 6486 823 0 otrip_decoded[4]
rlabel metal2 7774 1520 7774 1520 0 otrip_decoded[5]
rlabel metal2 7130 1656 7130 1656 0 otrip_decoded[6]
rlabel metal2 8418 1520 8418 1520 0 otrip_decoded[7]
rlabel metal2 9614 6749 9614 6749 0 outb_unbuf
rlabel metal2 9614 8279 9614 8279 0 timed_out
rlabel metal1 8188 10642 8188 10642 0 vtrip[0]
rlabel metal1 1886 10642 1886 10642 0 vtrip[1]
rlabel metal1 2668 10642 2668 10642 0 vtrip[2]
rlabel metal1 5336 10778 5336 10778 0 vtrip_decoded[0]
rlabel metal1 4048 10778 4048 10778 0 vtrip_decoded[1]
rlabel metal2 3266 11400 3266 11400 0 vtrip_decoded[2]
rlabel metal1 7912 10234 7912 10234 0 vtrip_decoded[3]
rlabel metal1 4692 10778 4692 10778 0 vtrip_decoded[4]
rlabel metal1 6624 10778 6624 10778 0 vtrip_decoded[5]
rlabel metal1 5888 10778 5888 10778 0 vtrip_decoded[6]
rlabel metal1 7222 10778 7222 10778 0 vtrip_decoded[7]
<< properties >>
string FIXED_BBOX 0 0 11173 13317
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712352531
<< nwell >>
rect -6235 -797 6235 797
<< mvpmos >>
rect -5977 -500 -5177 500
rect -5119 -500 -4319 500
rect -4261 -500 -3461 500
rect -3403 -500 -2603 500
rect -2545 -500 -1745 500
rect -1687 -500 -887 500
rect -829 -500 -29 500
rect 29 -500 829 500
rect 887 -500 1687 500
rect 1745 -500 2545 500
rect 2603 -500 3403 500
rect 3461 -500 4261 500
rect 4319 -500 5119 500
rect 5177 -500 5977 500
<< mvpdiff >>
rect -6035 488 -5977 500
rect -6035 -488 -6023 488
rect -5989 -488 -5977 488
rect -6035 -500 -5977 -488
rect -5177 488 -5119 500
rect -5177 -488 -5165 488
rect -5131 -488 -5119 488
rect -5177 -500 -5119 -488
rect -4319 488 -4261 500
rect -4319 -488 -4307 488
rect -4273 -488 -4261 488
rect -4319 -500 -4261 -488
rect -3461 488 -3403 500
rect -3461 -488 -3449 488
rect -3415 -488 -3403 488
rect -3461 -500 -3403 -488
rect -2603 488 -2545 500
rect -2603 -488 -2591 488
rect -2557 -488 -2545 488
rect -2603 -500 -2545 -488
rect -1745 488 -1687 500
rect -1745 -488 -1733 488
rect -1699 -488 -1687 488
rect -1745 -500 -1687 -488
rect -887 488 -829 500
rect -887 -488 -875 488
rect -841 -488 -829 488
rect -887 -500 -829 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 829 488 887 500
rect 829 -488 841 488
rect 875 -488 887 488
rect 829 -500 887 -488
rect 1687 488 1745 500
rect 1687 -488 1699 488
rect 1733 -488 1745 488
rect 1687 -500 1745 -488
rect 2545 488 2603 500
rect 2545 -488 2557 488
rect 2591 -488 2603 488
rect 2545 -500 2603 -488
rect 3403 488 3461 500
rect 3403 -488 3415 488
rect 3449 -488 3461 488
rect 3403 -500 3461 -488
rect 4261 488 4319 500
rect 4261 -488 4273 488
rect 4307 -488 4319 488
rect 4261 -500 4319 -488
rect 5119 488 5177 500
rect 5119 -488 5131 488
rect 5165 -488 5177 488
rect 5119 -500 5177 -488
rect 5977 488 6035 500
rect 5977 -488 5989 488
rect 6023 -488 6035 488
rect 5977 -500 6035 -488
<< mvpdiffc >>
rect -6023 -488 -5989 488
rect -5165 -488 -5131 488
rect -4307 -488 -4273 488
rect -3449 -488 -3415 488
rect -2591 -488 -2557 488
rect -1733 -488 -1699 488
rect -875 -488 -841 488
rect -17 -488 17 488
rect 841 -488 875 488
rect 1699 -488 1733 488
rect 2557 -488 2591 488
rect 3415 -488 3449 488
rect 4273 -488 4307 488
rect 5131 -488 5165 488
rect 5989 -488 6023 488
<< mvnsubdiff >>
rect -6169 719 6169 731
rect -6169 685 -6061 719
rect 6061 685 6169 719
rect -6169 673 6169 685
rect -6169 623 -6111 673
rect -6169 -623 -6157 623
rect -6123 -623 -6111 623
rect 6111 623 6169 673
rect -6169 -673 -6111 -623
rect 6111 -623 6123 623
rect 6157 -623 6169 623
rect 6111 -673 6169 -623
rect -6169 -685 6169 -673
rect -6169 -719 -6061 -685
rect 6061 -719 6169 -685
rect -6169 -731 6169 -719
<< mvnsubdiffcont >>
rect -6061 685 6061 719
rect -6157 -623 -6123 623
rect 6123 -623 6157 623
rect -6061 -719 6061 -685
<< poly >>
rect -5977 581 -5177 597
rect -5977 547 -5961 581
rect -5193 547 -5177 581
rect -5977 500 -5177 547
rect -5119 581 -4319 597
rect -5119 547 -5103 581
rect -4335 547 -4319 581
rect -5119 500 -4319 547
rect -4261 581 -3461 597
rect -4261 547 -4245 581
rect -3477 547 -3461 581
rect -4261 500 -3461 547
rect -3403 581 -2603 597
rect -3403 547 -3387 581
rect -2619 547 -2603 581
rect -3403 500 -2603 547
rect -2545 581 -1745 597
rect -2545 547 -2529 581
rect -1761 547 -1745 581
rect -2545 500 -1745 547
rect -1687 581 -887 597
rect -1687 547 -1671 581
rect -903 547 -887 581
rect -1687 500 -887 547
rect -829 581 -29 597
rect -829 547 -813 581
rect -45 547 -29 581
rect -829 500 -29 547
rect 29 581 829 597
rect 29 547 45 581
rect 813 547 829 581
rect 29 500 829 547
rect 887 581 1687 597
rect 887 547 903 581
rect 1671 547 1687 581
rect 887 500 1687 547
rect 1745 581 2545 597
rect 1745 547 1761 581
rect 2529 547 2545 581
rect 1745 500 2545 547
rect 2603 581 3403 597
rect 2603 547 2619 581
rect 3387 547 3403 581
rect 2603 500 3403 547
rect 3461 581 4261 597
rect 3461 547 3477 581
rect 4245 547 4261 581
rect 3461 500 4261 547
rect 4319 581 5119 597
rect 4319 547 4335 581
rect 5103 547 5119 581
rect 4319 500 5119 547
rect 5177 581 5977 597
rect 5177 547 5193 581
rect 5961 547 5977 581
rect 5177 500 5977 547
rect -5977 -547 -5177 -500
rect -5977 -581 -5961 -547
rect -5193 -581 -5177 -547
rect -5977 -597 -5177 -581
rect -5119 -547 -4319 -500
rect -5119 -581 -5103 -547
rect -4335 -581 -4319 -547
rect -5119 -597 -4319 -581
rect -4261 -547 -3461 -500
rect -4261 -581 -4245 -547
rect -3477 -581 -3461 -547
rect -4261 -597 -3461 -581
rect -3403 -547 -2603 -500
rect -3403 -581 -3387 -547
rect -2619 -581 -2603 -547
rect -3403 -597 -2603 -581
rect -2545 -547 -1745 -500
rect -2545 -581 -2529 -547
rect -1761 -581 -1745 -547
rect -2545 -597 -1745 -581
rect -1687 -547 -887 -500
rect -1687 -581 -1671 -547
rect -903 -581 -887 -547
rect -1687 -597 -887 -581
rect -829 -547 -29 -500
rect -829 -581 -813 -547
rect -45 -581 -29 -547
rect -829 -597 -29 -581
rect 29 -547 829 -500
rect 29 -581 45 -547
rect 813 -581 829 -547
rect 29 -597 829 -581
rect 887 -547 1687 -500
rect 887 -581 903 -547
rect 1671 -581 1687 -547
rect 887 -597 1687 -581
rect 1745 -547 2545 -500
rect 1745 -581 1761 -547
rect 2529 -581 2545 -547
rect 1745 -597 2545 -581
rect 2603 -547 3403 -500
rect 2603 -581 2619 -547
rect 3387 -581 3403 -547
rect 2603 -597 3403 -581
rect 3461 -547 4261 -500
rect 3461 -581 3477 -547
rect 4245 -581 4261 -547
rect 3461 -597 4261 -581
rect 4319 -547 5119 -500
rect 4319 -581 4335 -547
rect 5103 -581 5119 -547
rect 4319 -597 5119 -581
rect 5177 -547 5977 -500
rect 5177 -581 5193 -547
rect 5961 -581 5977 -547
rect 5177 -597 5977 -581
<< polycont >>
rect -5961 547 -5193 581
rect -5103 547 -4335 581
rect -4245 547 -3477 581
rect -3387 547 -2619 581
rect -2529 547 -1761 581
rect -1671 547 -903 581
rect -813 547 -45 581
rect 45 547 813 581
rect 903 547 1671 581
rect 1761 547 2529 581
rect 2619 547 3387 581
rect 3477 547 4245 581
rect 4335 547 5103 581
rect 5193 547 5961 581
rect -5961 -581 -5193 -547
rect -5103 -581 -4335 -547
rect -4245 -581 -3477 -547
rect -3387 -581 -2619 -547
rect -2529 -581 -1761 -547
rect -1671 -581 -903 -547
rect -813 -581 -45 -547
rect 45 -581 813 -547
rect 903 -581 1671 -547
rect 1761 -581 2529 -547
rect 2619 -581 3387 -547
rect 3477 -581 4245 -547
rect 4335 -581 5103 -547
rect 5193 -581 5961 -547
<< locali >>
rect -6157 685 -6061 719
rect 6061 685 6157 719
rect -6157 623 -6123 685
rect 6123 623 6157 685
rect -5977 547 -5961 581
rect -5193 547 -5177 581
rect -5119 547 -5103 581
rect -4335 547 -4319 581
rect -4261 547 -4245 581
rect -3477 547 -3461 581
rect -3403 547 -3387 581
rect -2619 547 -2603 581
rect -2545 547 -2529 581
rect -1761 547 -1745 581
rect -1687 547 -1671 581
rect -903 547 -887 581
rect -829 547 -813 581
rect -45 547 -29 581
rect 29 547 45 581
rect 813 547 829 581
rect 887 547 903 581
rect 1671 547 1687 581
rect 1745 547 1761 581
rect 2529 547 2545 581
rect 2603 547 2619 581
rect 3387 547 3403 581
rect 3461 547 3477 581
rect 4245 547 4261 581
rect 4319 547 4335 581
rect 5103 547 5119 581
rect 5177 547 5193 581
rect 5961 547 5977 581
rect -6023 488 -5989 504
rect -6023 -504 -5989 -488
rect -5165 488 -5131 504
rect -5165 -504 -5131 -488
rect -4307 488 -4273 504
rect -4307 -504 -4273 -488
rect -3449 488 -3415 504
rect -3449 -504 -3415 -488
rect -2591 488 -2557 504
rect -2591 -504 -2557 -488
rect -1733 488 -1699 504
rect -1733 -504 -1699 -488
rect -875 488 -841 504
rect -875 -504 -841 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 841 488 875 504
rect 841 -504 875 -488
rect 1699 488 1733 504
rect 1699 -504 1733 -488
rect 2557 488 2591 504
rect 2557 -504 2591 -488
rect 3415 488 3449 504
rect 3415 -504 3449 -488
rect 4273 488 4307 504
rect 4273 -504 4307 -488
rect 5131 488 5165 504
rect 5131 -504 5165 -488
rect 5989 488 6023 504
rect 5989 -504 6023 -488
rect -5977 -581 -5961 -547
rect -5193 -581 -5177 -547
rect -5119 -581 -5103 -547
rect -4335 -581 -4319 -547
rect -4261 -581 -4245 -547
rect -3477 -581 -3461 -547
rect -3403 -581 -3387 -547
rect -2619 -581 -2603 -547
rect -2545 -581 -2529 -547
rect -1761 -581 -1745 -547
rect -1687 -581 -1671 -547
rect -903 -581 -887 -547
rect -829 -581 -813 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 813 -581 829 -547
rect 887 -581 903 -547
rect 1671 -581 1687 -547
rect 1745 -581 1761 -547
rect 2529 -581 2545 -547
rect 2603 -581 2619 -547
rect 3387 -581 3403 -547
rect 3461 -581 3477 -547
rect 4245 -581 4261 -547
rect 4319 -581 4335 -547
rect 5103 -581 5119 -547
rect 5177 -581 5193 -547
rect 5961 -581 5977 -547
rect -6157 -685 -6123 -623
rect 6123 -685 6157 -623
rect -6157 -719 -6061 -685
rect 6061 -719 6157 -685
<< viali >>
rect -5961 547 -5193 581
rect -5103 547 -4335 581
rect -4245 547 -3477 581
rect -3387 547 -2619 581
rect -2529 547 -1761 581
rect -1671 547 -903 581
rect -813 547 -45 581
rect 45 547 813 581
rect 903 547 1671 581
rect 1761 547 2529 581
rect 2619 547 3387 581
rect 3477 547 4245 581
rect 4335 547 5103 581
rect 5193 547 5961 581
rect -6023 -488 -5989 488
rect -5165 -488 -5131 488
rect -4307 -488 -4273 488
rect -3449 -488 -3415 488
rect -2591 -488 -2557 488
rect -1733 -488 -1699 488
rect -875 -488 -841 488
rect -17 -488 17 488
rect 841 -488 875 488
rect 1699 -488 1733 488
rect 2557 -488 2591 488
rect 3415 -488 3449 488
rect 4273 -488 4307 488
rect 5131 -488 5165 488
rect 5989 -488 6023 488
rect -5961 -581 -5193 -547
rect -5103 -581 -4335 -547
rect -4245 -581 -3477 -547
rect -3387 -581 -2619 -547
rect -2529 -581 -1761 -547
rect -1671 -581 -903 -547
rect -813 -581 -45 -547
rect 45 -581 813 -547
rect 903 -581 1671 -547
rect 1761 -581 2529 -547
rect 2619 -581 3387 -547
rect 3477 -581 4245 -547
rect 4335 -581 5103 -547
rect 5193 -581 5961 -547
<< metal1 >>
rect -5973 581 -5181 587
rect -5973 547 -5961 581
rect -5193 547 -5181 581
rect -5973 541 -5181 547
rect -5115 581 -4323 587
rect -5115 547 -5103 581
rect -4335 547 -4323 581
rect -5115 541 -4323 547
rect -4257 581 -3465 587
rect -4257 547 -4245 581
rect -3477 547 -3465 581
rect -4257 541 -3465 547
rect -3399 581 -2607 587
rect -3399 547 -3387 581
rect -2619 547 -2607 581
rect -3399 541 -2607 547
rect -2541 581 -1749 587
rect -2541 547 -2529 581
rect -1761 547 -1749 581
rect -2541 541 -1749 547
rect -1683 581 -891 587
rect -1683 547 -1671 581
rect -903 547 -891 581
rect -1683 541 -891 547
rect -825 581 -33 587
rect -825 547 -813 581
rect -45 547 -33 581
rect -825 541 -33 547
rect 33 581 825 587
rect 33 547 45 581
rect 813 547 825 581
rect 33 541 825 547
rect 891 581 1683 587
rect 891 547 903 581
rect 1671 547 1683 581
rect 891 541 1683 547
rect 1749 581 2541 587
rect 1749 547 1761 581
rect 2529 547 2541 581
rect 1749 541 2541 547
rect 2607 581 3399 587
rect 2607 547 2619 581
rect 3387 547 3399 581
rect 2607 541 3399 547
rect 3465 581 4257 587
rect 3465 547 3477 581
rect 4245 547 4257 581
rect 3465 541 4257 547
rect 4323 581 5115 587
rect 4323 547 4335 581
rect 5103 547 5115 581
rect 4323 541 5115 547
rect 5181 581 5973 587
rect 5181 547 5193 581
rect 5961 547 5973 581
rect 5181 541 5973 547
rect -6029 488 -5983 500
rect -6029 -488 -6023 488
rect -5989 -488 -5983 488
rect -6029 -500 -5983 -488
rect -5171 488 -5125 500
rect -5171 -488 -5165 488
rect -5131 -488 -5125 488
rect -5171 -500 -5125 -488
rect -4313 488 -4267 500
rect -4313 -488 -4307 488
rect -4273 -488 -4267 488
rect -4313 -500 -4267 -488
rect -3455 488 -3409 500
rect -3455 -488 -3449 488
rect -3415 -488 -3409 488
rect -3455 -500 -3409 -488
rect -2597 488 -2551 500
rect -2597 -488 -2591 488
rect -2557 -488 -2551 488
rect -2597 -500 -2551 -488
rect -1739 488 -1693 500
rect -1739 -488 -1733 488
rect -1699 -488 -1693 488
rect -1739 -500 -1693 -488
rect -881 488 -835 500
rect -881 -488 -875 488
rect -841 -488 -835 488
rect -881 -500 -835 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 835 488 881 500
rect 835 -488 841 488
rect 875 -488 881 488
rect 835 -500 881 -488
rect 1693 488 1739 500
rect 1693 -488 1699 488
rect 1733 -488 1739 488
rect 1693 -500 1739 -488
rect 2551 488 2597 500
rect 2551 -488 2557 488
rect 2591 -488 2597 488
rect 2551 -500 2597 -488
rect 3409 488 3455 500
rect 3409 -488 3415 488
rect 3449 -488 3455 488
rect 3409 -500 3455 -488
rect 4267 488 4313 500
rect 4267 -488 4273 488
rect 4307 -488 4313 488
rect 4267 -500 4313 -488
rect 5125 488 5171 500
rect 5125 -488 5131 488
rect 5165 -488 5171 488
rect 5125 -500 5171 -488
rect 5983 488 6029 500
rect 5983 -488 5989 488
rect 6023 -488 6029 488
rect 5983 -500 6029 -488
rect -5973 -547 -5181 -541
rect -5973 -581 -5961 -547
rect -5193 -581 -5181 -547
rect -5973 -587 -5181 -581
rect -5115 -547 -4323 -541
rect -5115 -581 -5103 -547
rect -4335 -581 -4323 -547
rect -5115 -587 -4323 -581
rect -4257 -547 -3465 -541
rect -4257 -581 -4245 -547
rect -3477 -581 -3465 -547
rect -4257 -587 -3465 -581
rect -3399 -547 -2607 -541
rect -3399 -581 -3387 -547
rect -2619 -581 -2607 -547
rect -3399 -587 -2607 -581
rect -2541 -547 -1749 -541
rect -2541 -581 -2529 -547
rect -1761 -581 -1749 -547
rect -2541 -587 -1749 -581
rect -1683 -547 -891 -541
rect -1683 -581 -1671 -547
rect -903 -581 -891 -547
rect -1683 -587 -891 -581
rect -825 -547 -33 -541
rect -825 -581 -813 -547
rect -45 -581 -33 -547
rect -825 -587 -33 -581
rect 33 -547 825 -541
rect 33 -581 45 -547
rect 813 -581 825 -547
rect 33 -587 825 -581
rect 891 -547 1683 -541
rect 891 -581 903 -547
rect 1671 -581 1683 -547
rect 891 -587 1683 -581
rect 1749 -547 2541 -541
rect 1749 -581 1761 -547
rect 2529 -581 2541 -547
rect 1749 -587 2541 -581
rect 2607 -547 3399 -541
rect 2607 -581 2619 -547
rect 3387 -581 3399 -547
rect 2607 -587 3399 -581
rect 3465 -547 4257 -541
rect 3465 -581 3477 -547
rect 4245 -581 4257 -547
rect 3465 -587 4257 -581
rect 4323 -547 5115 -541
rect 4323 -581 4335 -547
rect 5103 -581 5115 -547
rect 4323 -587 5115 -581
rect 5181 -547 5973 -541
rect 5181 -581 5193 -547
rect 5961 -581 5973 -547
rect 5181 -587 5973 -581
<< properties >>
string FIXED_BBOX -6140 -702 6140 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 4 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

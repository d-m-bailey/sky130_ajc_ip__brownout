magic
tech sky130A
magscale 1 2
timestamp 1712722749
<< nwell >>
rect -618 -164 618 198
<< pmos >>
rect -524 -64 -424 136
rect -366 -64 -266 136
rect -208 -64 -108 136
rect -50 -64 50 136
rect 108 -64 208 136
rect 266 -64 366 136
rect 424 -64 524 136
<< pdiff >>
rect -582 124 -524 136
rect -582 -52 -570 124
rect -536 -52 -524 124
rect -582 -64 -524 -52
rect -424 124 -366 136
rect -424 -52 -412 124
rect -378 -52 -366 124
rect -424 -64 -366 -52
rect -266 124 -208 136
rect -266 -52 -254 124
rect -220 -52 -208 124
rect -266 -64 -208 -52
rect -108 124 -50 136
rect -108 -52 -96 124
rect -62 -52 -50 124
rect -108 -64 -50 -52
rect 50 124 108 136
rect 50 -52 62 124
rect 96 -52 108 124
rect 50 -64 108 -52
rect 208 124 266 136
rect 208 -52 220 124
rect 254 -52 266 124
rect 208 -64 266 -52
rect 366 124 424 136
rect 366 -52 378 124
rect 412 -52 424 124
rect 366 -64 424 -52
rect 524 124 582 136
rect 524 -52 536 124
rect 570 -52 582 124
rect 524 -64 582 -52
<< pdiffc >>
rect -570 -52 -536 124
rect -412 -52 -378 124
rect -254 -52 -220 124
rect -96 -52 -62 124
rect 62 -52 96 124
rect 220 -52 254 124
rect 378 -52 412 124
rect 536 -52 570 124
<< poly >>
rect -524 136 -424 162
rect -366 136 -266 162
rect -208 136 -108 162
rect -50 136 50 162
rect 108 136 208 162
rect 266 136 366 162
rect 424 136 524 162
rect -524 -111 -424 -64
rect -524 -145 -508 -111
rect -440 -145 -424 -111
rect -524 -161 -424 -145
rect -366 -111 -266 -64
rect -366 -145 -350 -111
rect -282 -145 -266 -111
rect -366 -161 -266 -145
rect -208 -111 -108 -64
rect -208 -145 -192 -111
rect -124 -145 -108 -111
rect -208 -161 -108 -145
rect -50 -111 50 -64
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect -50 -161 50 -145
rect 108 -111 208 -64
rect 108 -145 124 -111
rect 192 -145 208 -111
rect 108 -161 208 -145
rect 266 -111 366 -64
rect 266 -145 282 -111
rect 350 -145 366 -111
rect 266 -161 366 -145
rect 424 -111 524 -64
rect 424 -145 440 -111
rect 508 -145 524 -111
rect 424 -161 524 -145
<< polycont >>
rect -508 -145 -440 -111
rect -350 -145 -282 -111
rect -192 -145 -124 -111
rect -34 -145 34 -111
rect 124 -145 192 -111
rect 282 -145 350 -111
rect 440 -145 508 -111
<< locali >>
rect -570 124 -536 140
rect -570 -68 -536 -52
rect -412 124 -378 140
rect -412 -68 -378 -52
rect -254 124 -220 140
rect -254 -68 -220 -52
rect -96 124 -62 140
rect -96 -68 -62 -52
rect 62 124 96 140
rect 62 -68 96 -52
rect 220 124 254 140
rect 220 -68 254 -52
rect 378 124 412 140
rect 378 -68 412 -52
rect 536 124 570 140
rect 536 -68 570 -52
rect -524 -145 -508 -111
rect -440 -145 -424 -111
rect -366 -145 -350 -111
rect -282 -145 -266 -111
rect -208 -145 -192 -111
rect -124 -145 -108 -111
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect 108 -145 124 -111
rect 192 -145 208 -111
rect 266 -145 282 -111
rect 350 -145 366 -111
rect 424 -145 440 -111
rect 508 -145 524 -111
<< viali >>
rect -570 -52 -536 124
rect -412 -52 -378 124
rect -254 -52 -220 124
rect -96 -52 -62 124
rect 62 -52 96 124
rect 220 -52 254 124
rect 378 -52 412 124
rect 536 -52 570 124
rect -508 -145 -440 -111
rect -350 -145 -282 -111
rect -192 -145 -124 -111
rect -34 -145 34 -111
rect 124 -145 192 -111
rect 282 -145 350 -111
rect 440 -145 508 -111
<< metal1 >>
rect -576 124 -530 136
rect -576 -52 -570 124
rect -536 -52 -530 124
rect -576 -64 -530 -52
rect -418 124 -372 136
rect -418 -52 -412 124
rect -378 -52 -372 124
rect -418 -64 -372 -52
rect -260 124 -214 136
rect -260 -52 -254 124
rect -220 -52 -214 124
rect -260 -64 -214 -52
rect -102 124 -56 136
rect -102 -52 -96 124
rect -62 -52 -56 124
rect -102 -64 -56 -52
rect 56 124 102 136
rect 56 -52 62 124
rect 96 -52 102 124
rect 56 -64 102 -52
rect 214 124 260 136
rect 214 -52 220 124
rect 254 -52 260 124
rect 214 -64 260 -52
rect 372 124 418 136
rect 372 -52 378 124
rect 412 -52 418 124
rect 372 -64 418 -52
rect 530 124 576 136
rect 530 -52 536 124
rect 570 -52 576 124
rect 530 -64 576 -52
rect -520 -111 -428 -105
rect -520 -145 -508 -111
rect -440 -145 -428 -111
rect -520 -151 -428 -145
rect -362 -111 -270 -105
rect -362 -145 -350 -111
rect -282 -145 -270 -111
rect -362 -151 -270 -145
rect -204 -111 -112 -105
rect -204 -145 -192 -111
rect -124 -145 -112 -111
rect -204 -151 -112 -145
rect -46 -111 46 -105
rect -46 -145 -34 -111
rect 34 -145 46 -111
rect -46 -151 46 -145
rect 112 -111 204 -105
rect 112 -145 124 -111
rect 192 -145 204 -111
rect 112 -151 204 -145
rect 270 -111 362 -105
rect 270 -145 282 -111
rect 350 -145 362 -111
rect 270 -151 362 -145
rect 428 -111 520 -105
rect 428 -145 440 -111
rect 508 -145 520 -111
rect 428 -151 520 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 7 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712709231
<< pwell >>
rect -2197 -10082 2197 10082
<< psubdiff >>
rect -2161 10012 -2065 10046
rect 2065 10012 2161 10046
rect -2161 9950 -2127 10012
rect 2127 9950 2161 10012
rect -2161 -10012 -2127 -9950
rect 2127 -10012 2161 -9950
rect -2161 -10046 -2065 -10012
rect 2065 -10046 2161 -10012
<< psubdiffcont >>
rect -2065 10012 2065 10046
rect -2161 -9950 -2127 9950
rect 2127 -9950 2161 9950
rect -2065 -10046 2065 -10012
<< xpolycontact >>
rect -2031 9484 -1749 9916
rect -2031 -9916 -1749 -9484
rect -1653 9484 -1371 9916
rect -1653 -9916 -1371 -9484
rect -1275 9484 -993 9916
rect -1275 -9916 -993 -9484
rect -897 9484 -615 9916
rect -897 -9916 -615 -9484
rect -519 9484 -237 9916
rect -519 -9916 -237 -9484
rect -141 9484 141 9916
rect -141 -9916 141 -9484
rect 237 9484 519 9916
rect 237 -9916 519 -9484
rect 615 9484 897 9916
rect 615 -9916 897 -9484
rect 993 9484 1275 9916
rect 993 -9916 1275 -9484
rect 1371 9484 1653 9916
rect 1371 -9916 1653 -9484
rect 1749 9484 2031 9916
rect 1749 -9916 2031 -9484
<< xpolyres >>
rect -2031 -9484 -1749 9484
rect -1653 -9484 -1371 9484
rect -1275 -9484 -993 9484
rect -897 -9484 -615 9484
rect -519 -9484 -237 9484
rect -141 -9484 141 9484
rect 237 -9484 519 9484
rect 615 -9484 897 9484
rect 993 -9484 1275 9484
rect 1371 -9484 1653 9484
rect 1749 -9484 2031 9484
<< locali >>
rect -2161 10012 -2065 10046
rect 2065 10012 2161 10046
rect -2161 9950 -2127 10012
rect 2127 9950 2161 10012
rect -2161 -10012 -2127 -9950
rect 2127 -10012 2161 -9950
rect -2161 -10046 -2065 -10012
rect 2065 -10046 2161 -10012
<< viali >>
rect -2015 9501 -1765 9898
rect -1637 9501 -1387 9898
rect -1259 9501 -1009 9898
rect -881 9501 -631 9898
rect -503 9501 -253 9898
rect -125 9501 125 9898
rect 253 9501 503 9898
rect 631 9501 881 9898
rect 1009 9501 1259 9898
rect 1387 9501 1637 9898
rect 1765 9501 2015 9898
rect -2015 -9898 -1765 -9501
rect -1637 -9898 -1387 -9501
rect -1259 -9898 -1009 -9501
rect -881 -9898 -631 -9501
rect -503 -9898 -253 -9501
rect -125 -9898 125 -9501
rect 253 -9898 503 -9501
rect 631 -9898 881 -9501
rect 1009 -9898 1259 -9501
rect 1387 -9898 1637 -9501
rect 1765 -9898 2015 -9501
<< metal1 >>
rect -2021 9898 -1759 9910
rect -2021 9501 -2015 9898
rect -1765 9501 -1759 9898
rect -2021 9489 -1759 9501
rect -1643 9898 -1381 9910
rect -1643 9501 -1637 9898
rect -1387 9501 -1381 9898
rect -1643 9489 -1381 9501
rect -1265 9898 -1003 9910
rect -1265 9501 -1259 9898
rect -1009 9501 -1003 9898
rect -1265 9489 -1003 9501
rect -887 9898 -625 9910
rect -887 9501 -881 9898
rect -631 9501 -625 9898
rect -887 9489 -625 9501
rect -509 9898 -247 9910
rect -509 9501 -503 9898
rect -253 9501 -247 9898
rect -509 9489 -247 9501
rect -131 9898 131 9910
rect -131 9501 -125 9898
rect 125 9501 131 9898
rect -131 9489 131 9501
rect 247 9898 509 9910
rect 247 9501 253 9898
rect 503 9501 509 9898
rect 247 9489 509 9501
rect 625 9898 887 9910
rect 625 9501 631 9898
rect 881 9501 887 9898
rect 625 9489 887 9501
rect 1003 9898 1265 9910
rect 1003 9501 1009 9898
rect 1259 9501 1265 9898
rect 1003 9489 1265 9501
rect 1381 9898 1643 9910
rect 1381 9501 1387 9898
rect 1637 9501 1643 9898
rect 1381 9489 1643 9501
rect 1759 9898 2021 9910
rect 1759 9501 1765 9898
rect 2015 9501 2021 9898
rect 1759 9489 2021 9501
rect -2021 -9501 -1759 -9489
rect -2021 -9898 -2015 -9501
rect -1765 -9898 -1759 -9501
rect -2021 -9910 -1759 -9898
rect -1643 -9501 -1381 -9489
rect -1643 -9898 -1637 -9501
rect -1387 -9898 -1381 -9501
rect -1643 -9910 -1381 -9898
rect -1265 -9501 -1003 -9489
rect -1265 -9898 -1259 -9501
rect -1009 -9898 -1003 -9501
rect -1265 -9910 -1003 -9898
rect -887 -9501 -625 -9489
rect -887 -9898 -881 -9501
rect -631 -9898 -625 -9501
rect -887 -9910 -625 -9898
rect -509 -9501 -247 -9489
rect -509 -9898 -503 -9501
rect -253 -9898 -247 -9501
rect -509 -9910 -247 -9898
rect -131 -9501 131 -9489
rect -131 -9898 -125 -9501
rect 125 -9898 131 -9501
rect -131 -9910 131 -9898
rect 247 -9501 509 -9489
rect 247 -9898 253 -9501
rect 503 -9898 509 -9501
rect 247 -9910 509 -9898
rect 625 -9501 887 -9489
rect 625 -9898 631 -9501
rect 881 -9898 887 -9501
rect 625 -9910 887 -9898
rect 1003 -9501 1265 -9489
rect 1003 -9898 1009 -9501
rect 1259 -9898 1265 -9501
rect 1003 -9910 1265 -9898
rect 1381 -9501 1643 -9489
rect 1381 -9898 1387 -9501
rect 1637 -9898 1643 -9501
rect 1381 -9910 1643 -9898
rect 1759 -9501 2021 -9489
rect 1759 -9898 1765 -9501
rect 2015 -9898 2021 -9501
rect 1759 -9910 2021 -9898
<< properties >>
string FIXED_BBOX -2144 -10029 2144 10029
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 95 m 1 nx 11 wmin 1.410 lmin 0.50 rho 2000 val 135.018k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712594819
<< pwell >>
rect -13348 -4082 13348 4082
<< psubdiff >>
rect -13312 4012 -13216 4046
rect 13216 4012 13312 4046
rect -13312 3950 -13278 4012
rect 13278 3950 13312 4012
rect -13312 -4012 -13278 -3950
rect 13278 -4012 13312 -3950
rect -13312 -4046 -13216 -4012
rect 13216 -4046 13312 -4012
<< psubdiffcont >>
rect -13216 4012 13216 4046
rect -13312 -3950 -13278 3950
rect 13278 -3950 13312 3950
rect -13216 -4046 13216 -4012
<< xpolycontact >>
rect -13182 3484 -12900 3916
rect -13182 -3916 -12900 -3484
rect -12804 3484 -12522 3916
rect -12804 -3916 -12522 -3484
rect -12426 3484 -12144 3916
rect -12426 -3916 -12144 -3484
rect -12048 3484 -11766 3916
rect -12048 -3916 -11766 -3484
rect -11670 3484 -11388 3916
rect -11670 -3916 -11388 -3484
rect -11292 3484 -11010 3916
rect -11292 -3916 -11010 -3484
rect -10914 3484 -10632 3916
rect -10914 -3916 -10632 -3484
rect -10536 3484 -10254 3916
rect -10536 -3916 -10254 -3484
rect -10158 3484 -9876 3916
rect -10158 -3916 -9876 -3484
rect -9780 3484 -9498 3916
rect -9780 -3916 -9498 -3484
rect -9402 3484 -9120 3916
rect -9402 -3916 -9120 -3484
rect -9024 3484 -8742 3916
rect -9024 -3916 -8742 -3484
rect -8646 3484 -8364 3916
rect -8646 -3916 -8364 -3484
rect -8268 3484 -7986 3916
rect -8268 -3916 -7986 -3484
rect -7890 3484 -7608 3916
rect -7890 -3916 -7608 -3484
rect -7512 3484 -7230 3916
rect -7512 -3916 -7230 -3484
rect -7134 3484 -6852 3916
rect -7134 -3916 -6852 -3484
rect -6756 3484 -6474 3916
rect -6756 -3916 -6474 -3484
rect -6378 3484 -6096 3916
rect -6378 -3916 -6096 -3484
rect -6000 3484 -5718 3916
rect -6000 -3916 -5718 -3484
rect -5622 3484 -5340 3916
rect -5622 -3916 -5340 -3484
rect -5244 3484 -4962 3916
rect -5244 -3916 -4962 -3484
rect -4866 3484 -4584 3916
rect -4866 -3916 -4584 -3484
rect -4488 3484 -4206 3916
rect -4488 -3916 -4206 -3484
rect -4110 3484 -3828 3916
rect -4110 -3916 -3828 -3484
rect -3732 3484 -3450 3916
rect -3732 -3916 -3450 -3484
rect -3354 3484 -3072 3916
rect -3354 -3916 -3072 -3484
rect -2976 3484 -2694 3916
rect -2976 -3916 -2694 -3484
rect -2598 3484 -2316 3916
rect -2598 -3916 -2316 -3484
rect -2220 3484 -1938 3916
rect -2220 -3916 -1938 -3484
rect -1842 3484 -1560 3916
rect -1842 -3916 -1560 -3484
rect -1464 3484 -1182 3916
rect -1464 -3916 -1182 -3484
rect -1086 3484 -804 3916
rect -1086 -3916 -804 -3484
rect -708 3484 -426 3916
rect -708 -3916 -426 -3484
rect -330 3484 -48 3916
rect -330 -3916 -48 -3484
rect 48 3484 330 3916
rect 48 -3916 330 -3484
rect 426 3484 708 3916
rect 426 -3916 708 -3484
rect 804 3484 1086 3916
rect 804 -3916 1086 -3484
rect 1182 3484 1464 3916
rect 1182 -3916 1464 -3484
rect 1560 3484 1842 3916
rect 1560 -3916 1842 -3484
rect 1938 3484 2220 3916
rect 1938 -3916 2220 -3484
rect 2316 3484 2598 3916
rect 2316 -3916 2598 -3484
rect 2694 3484 2976 3916
rect 2694 -3916 2976 -3484
rect 3072 3484 3354 3916
rect 3072 -3916 3354 -3484
rect 3450 3484 3732 3916
rect 3450 -3916 3732 -3484
rect 3828 3484 4110 3916
rect 3828 -3916 4110 -3484
rect 4206 3484 4488 3916
rect 4206 -3916 4488 -3484
rect 4584 3484 4866 3916
rect 4584 -3916 4866 -3484
rect 4962 3484 5244 3916
rect 4962 -3916 5244 -3484
rect 5340 3484 5622 3916
rect 5340 -3916 5622 -3484
rect 5718 3484 6000 3916
rect 5718 -3916 6000 -3484
rect 6096 3484 6378 3916
rect 6096 -3916 6378 -3484
rect 6474 3484 6756 3916
rect 6474 -3916 6756 -3484
rect 6852 3484 7134 3916
rect 6852 -3916 7134 -3484
rect 7230 3484 7512 3916
rect 7230 -3916 7512 -3484
rect 7608 3484 7890 3916
rect 7608 -3916 7890 -3484
rect 7986 3484 8268 3916
rect 7986 -3916 8268 -3484
rect 8364 3484 8646 3916
rect 8364 -3916 8646 -3484
rect 8742 3484 9024 3916
rect 8742 -3916 9024 -3484
rect 9120 3484 9402 3916
rect 9120 -3916 9402 -3484
rect 9498 3484 9780 3916
rect 9498 -3916 9780 -3484
rect 9876 3484 10158 3916
rect 9876 -3916 10158 -3484
rect 10254 3484 10536 3916
rect 10254 -3916 10536 -3484
rect 10632 3484 10914 3916
rect 10632 -3916 10914 -3484
rect 11010 3484 11292 3916
rect 11010 -3916 11292 -3484
rect 11388 3484 11670 3916
rect 11388 -3916 11670 -3484
rect 11766 3484 12048 3916
rect 11766 -3916 12048 -3484
rect 12144 3484 12426 3916
rect 12144 -3916 12426 -3484
rect 12522 3484 12804 3916
rect 12522 -3916 12804 -3484
rect 12900 3484 13182 3916
rect 12900 -3916 13182 -3484
<< xpolyres >>
rect -13182 -3484 -12900 3484
rect -12804 -3484 -12522 3484
rect -12426 -3484 -12144 3484
rect -12048 -3484 -11766 3484
rect -11670 -3484 -11388 3484
rect -11292 -3484 -11010 3484
rect -10914 -3484 -10632 3484
rect -10536 -3484 -10254 3484
rect -10158 -3484 -9876 3484
rect -9780 -3484 -9498 3484
rect -9402 -3484 -9120 3484
rect -9024 -3484 -8742 3484
rect -8646 -3484 -8364 3484
rect -8268 -3484 -7986 3484
rect -7890 -3484 -7608 3484
rect -7512 -3484 -7230 3484
rect -7134 -3484 -6852 3484
rect -6756 -3484 -6474 3484
rect -6378 -3484 -6096 3484
rect -6000 -3484 -5718 3484
rect -5622 -3484 -5340 3484
rect -5244 -3484 -4962 3484
rect -4866 -3484 -4584 3484
rect -4488 -3484 -4206 3484
rect -4110 -3484 -3828 3484
rect -3732 -3484 -3450 3484
rect -3354 -3484 -3072 3484
rect -2976 -3484 -2694 3484
rect -2598 -3484 -2316 3484
rect -2220 -3484 -1938 3484
rect -1842 -3484 -1560 3484
rect -1464 -3484 -1182 3484
rect -1086 -3484 -804 3484
rect -708 -3484 -426 3484
rect -330 -3484 -48 3484
rect 48 -3484 330 3484
rect 426 -3484 708 3484
rect 804 -3484 1086 3484
rect 1182 -3484 1464 3484
rect 1560 -3484 1842 3484
rect 1938 -3484 2220 3484
rect 2316 -3484 2598 3484
rect 2694 -3484 2976 3484
rect 3072 -3484 3354 3484
rect 3450 -3484 3732 3484
rect 3828 -3484 4110 3484
rect 4206 -3484 4488 3484
rect 4584 -3484 4866 3484
rect 4962 -3484 5244 3484
rect 5340 -3484 5622 3484
rect 5718 -3484 6000 3484
rect 6096 -3484 6378 3484
rect 6474 -3484 6756 3484
rect 6852 -3484 7134 3484
rect 7230 -3484 7512 3484
rect 7608 -3484 7890 3484
rect 7986 -3484 8268 3484
rect 8364 -3484 8646 3484
rect 8742 -3484 9024 3484
rect 9120 -3484 9402 3484
rect 9498 -3484 9780 3484
rect 9876 -3484 10158 3484
rect 10254 -3484 10536 3484
rect 10632 -3484 10914 3484
rect 11010 -3484 11292 3484
rect 11388 -3484 11670 3484
rect 11766 -3484 12048 3484
rect 12144 -3484 12426 3484
rect 12522 -3484 12804 3484
rect 12900 -3484 13182 3484
<< locali >>
rect -13312 4012 -13216 4046
rect 13216 4012 13312 4046
rect -13312 3950 -13278 4012
rect 13278 3950 13312 4012
rect -13312 -4012 -13278 -3950
rect 13278 -4012 13312 -3950
rect -13312 -4046 -13216 -4012
rect 13216 -4046 13312 -4012
<< viali >>
rect -13166 3501 -12916 3898
rect -12788 3501 -12538 3898
rect -12410 3501 -12160 3898
rect -12032 3501 -11782 3898
rect -11654 3501 -11404 3898
rect -11276 3501 -11026 3898
rect -10898 3501 -10648 3898
rect -10520 3501 -10270 3898
rect -10142 3501 -9892 3898
rect -9764 3501 -9514 3898
rect -9386 3501 -9136 3898
rect -9008 3501 -8758 3898
rect -8630 3501 -8380 3898
rect -8252 3501 -8002 3898
rect -7874 3501 -7624 3898
rect -7496 3501 -7246 3898
rect -7118 3501 -6868 3898
rect -6740 3501 -6490 3898
rect -6362 3501 -6112 3898
rect -5984 3501 -5734 3898
rect -5606 3501 -5356 3898
rect -5228 3501 -4978 3898
rect -4850 3501 -4600 3898
rect -4472 3501 -4222 3898
rect -4094 3501 -3844 3898
rect -3716 3501 -3466 3898
rect -3338 3501 -3088 3898
rect -2960 3501 -2710 3898
rect -2582 3501 -2332 3898
rect -2204 3501 -1954 3898
rect -1826 3501 -1576 3898
rect -1448 3501 -1198 3898
rect -1070 3501 -820 3898
rect -692 3501 -442 3898
rect -314 3501 -64 3898
rect 64 3501 314 3898
rect 442 3501 692 3898
rect 820 3501 1070 3898
rect 1198 3501 1448 3898
rect 1576 3501 1826 3898
rect 1954 3501 2204 3898
rect 2332 3501 2582 3898
rect 2710 3501 2960 3898
rect 3088 3501 3338 3898
rect 3466 3501 3716 3898
rect 3844 3501 4094 3898
rect 4222 3501 4472 3898
rect 4600 3501 4850 3898
rect 4978 3501 5228 3898
rect 5356 3501 5606 3898
rect 5734 3501 5984 3898
rect 6112 3501 6362 3898
rect 6490 3501 6740 3898
rect 6868 3501 7118 3898
rect 7246 3501 7496 3898
rect 7624 3501 7874 3898
rect 8002 3501 8252 3898
rect 8380 3501 8630 3898
rect 8758 3501 9008 3898
rect 9136 3501 9386 3898
rect 9514 3501 9764 3898
rect 9892 3501 10142 3898
rect 10270 3501 10520 3898
rect 10648 3501 10898 3898
rect 11026 3501 11276 3898
rect 11404 3501 11654 3898
rect 11782 3501 12032 3898
rect 12160 3501 12410 3898
rect 12538 3501 12788 3898
rect 12916 3501 13166 3898
rect -13166 -3898 -12916 -3501
rect -12788 -3898 -12538 -3501
rect -12410 -3898 -12160 -3501
rect -12032 -3898 -11782 -3501
rect -11654 -3898 -11404 -3501
rect -11276 -3898 -11026 -3501
rect -10898 -3898 -10648 -3501
rect -10520 -3898 -10270 -3501
rect -10142 -3898 -9892 -3501
rect -9764 -3898 -9514 -3501
rect -9386 -3898 -9136 -3501
rect -9008 -3898 -8758 -3501
rect -8630 -3898 -8380 -3501
rect -8252 -3898 -8002 -3501
rect -7874 -3898 -7624 -3501
rect -7496 -3898 -7246 -3501
rect -7118 -3898 -6868 -3501
rect -6740 -3898 -6490 -3501
rect -6362 -3898 -6112 -3501
rect -5984 -3898 -5734 -3501
rect -5606 -3898 -5356 -3501
rect -5228 -3898 -4978 -3501
rect -4850 -3898 -4600 -3501
rect -4472 -3898 -4222 -3501
rect -4094 -3898 -3844 -3501
rect -3716 -3898 -3466 -3501
rect -3338 -3898 -3088 -3501
rect -2960 -3898 -2710 -3501
rect -2582 -3898 -2332 -3501
rect -2204 -3898 -1954 -3501
rect -1826 -3898 -1576 -3501
rect -1448 -3898 -1198 -3501
rect -1070 -3898 -820 -3501
rect -692 -3898 -442 -3501
rect -314 -3898 -64 -3501
rect 64 -3898 314 -3501
rect 442 -3898 692 -3501
rect 820 -3898 1070 -3501
rect 1198 -3898 1448 -3501
rect 1576 -3898 1826 -3501
rect 1954 -3898 2204 -3501
rect 2332 -3898 2582 -3501
rect 2710 -3898 2960 -3501
rect 3088 -3898 3338 -3501
rect 3466 -3898 3716 -3501
rect 3844 -3898 4094 -3501
rect 4222 -3898 4472 -3501
rect 4600 -3898 4850 -3501
rect 4978 -3898 5228 -3501
rect 5356 -3898 5606 -3501
rect 5734 -3898 5984 -3501
rect 6112 -3898 6362 -3501
rect 6490 -3898 6740 -3501
rect 6868 -3898 7118 -3501
rect 7246 -3898 7496 -3501
rect 7624 -3898 7874 -3501
rect 8002 -3898 8252 -3501
rect 8380 -3898 8630 -3501
rect 8758 -3898 9008 -3501
rect 9136 -3898 9386 -3501
rect 9514 -3898 9764 -3501
rect 9892 -3898 10142 -3501
rect 10270 -3898 10520 -3501
rect 10648 -3898 10898 -3501
rect 11026 -3898 11276 -3501
rect 11404 -3898 11654 -3501
rect 11782 -3898 12032 -3501
rect 12160 -3898 12410 -3501
rect 12538 -3898 12788 -3501
rect 12916 -3898 13166 -3501
<< metal1 >>
rect -13172 3898 -12910 3910
rect -13172 3501 -13166 3898
rect -12916 3501 -12910 3898
rect -13172 3489 -12910 3501
rect -12794 3898 -12532 3910
rect -12794 3501 -12788 3898
rect -12538 3501 -12532 3898
rect -12794 3489 -12532 3501
rect -12416 3898 -12154 3910
rect -12416 3501 -12410 3898
rect -12160 3501 -12154 3898
rect -12416 3489 -12154 3501
rect -12038 3898 -11776 3910
rect -12038 3501 -12032 3898
rect -11782 3501 -11776 3898
rect -12038 3489 -11776 3501
rect -11660 3898 -11398 3910
rect -11660 3501 -11654 3898
rect -11404 3501 -11398 3898
rect -11660 3489 -11398 3501
rect -11282 3898 -11020 3910
rect -11282 3501 -11276 3898
rect -11026 3501 -11020 3898
rect -11282 3489 -11020 3501
rect -10904 3898 -10642 3910
rect -10904 3501 -10898 3898
rect -10648 3501 -10642 3898
rect -10904 3489 -10642 3501
rect -10526 3898 -10264 3910
rect -10526 3501 -10520 3898
rect -10270 3501 -10264 3898
rect -10526 3489 -10264 3501
rect -10148 3898 -9886 3910
rect -10148 3501 -10142 3898
rect -9892 3501 -9886 3898
rect -10148 3489 -9886 3501
rect -9770 3898 -9508 3910
rect -9770 3501 -9764 3898
rect -9514 3501 -9508 3898
rect -9770 3489 -9508 3501
rect -9392 3898 -9130 3910
rect -9392 3501 -9386 3898
rect -9136 3501 -9130 3898
rect -9392 3489 -9130 3501
rect -9014 3898 -8752 3910
rect -9014 3501 -9008 3898
rect -8758 3501 -8752 3898
rect -9014 3489 -8752 3501
rect -8636 3898 -8374 3910
rect -8636 3501 -8630 3898
rect -8380 3501 -8374 3898
rect -8636 3489 -8374 3501
rect -8258 3898 -7996 3910
rect -8258 3501 -8252 3898
rect -8002 3501 -7996 3898
rect -8258 3489 -7996 3501
rect -7880 3898 -7618 3910
rect -7880 3501 -7874 3898
rect -7624 3501 -7618 3898
rect -7880 3489 -7618 3501
rect -7502 3898 -7240 3910
rect -7502 3501 -7496 3898
rect -7246 3501 -7240 3898
rect -7502 3489 -7240 3501
rect -7124 3898 -6862 3910
rect -7124 3501 -7118 3898
rect -6868 3501 -6862 3898
rect -7124 3489 -6862 3501
rect -6746 3898 -6484 3910
rect -6746 3501 -6740 3898
rect -6490 3501 -6484 3898
rect -6746 3489 -6484 3501
rect -6368 3898 -6106 3910
rect -6368 3501 -6362 3898
rect -6112 3501 -6106 3898
rect -6368 3489 -6106 3501
rect -5990 3898 -5728 3910
rect -5990 3501 -5984 3898
rect -5734 3501 -5728 3898
rect -5990 3489 -5728 3501
rect -5612 3898 -5350 3910
rect -5612 3501 -5606 3898
rect -5356 3501 -5350 3898
rect -5612 3489 -5350 3501
rect -5234 3898 -4972 3910
rect -5234 3501 -5228 3898
rect -4978 3501 -4972 3898
rect -5234 3489 -4972 3501
rect -4856 3898 -4594 3910
rect -4856 3501 -4850 3898
rect -4600 3501 -4594 3898
rect -4856 3489 -4594 3501
rect -4478 3898 -4216 3910
rect -4478 3501 -4472 3898
rect -4222 3501 -4216 3898
rect -4478 3489 -4216 3501
rect -4100 3898 -3838 3910
rect -4100 3501 -4094 3898
rect -3844 3501 -3838 3898
rect -4100 3489 -3838 3501
rect -3722 3898 -3460 3910
rect -3722 3501 -3716 3898
rect -3466 3501 -3460 3898
rect -3722 3489 -3460 3501
rect -3344 3898 -3082 3910
rect -3344 3501 -3338 3898
rect -3088 3501 -3082 3898
rect -3344 3489 -3082 3501
rect -2966 3898 -2704 3910
rect -2966 3501 -2960 3898
rect -2710 3501 -2704 3898
rect -2966 3489 -2704 3501
rect -2588 3898 -2326 3910
rect -2588 3501 -2582 3898
rect -2332 3501 -2326 3898
rect -2588 3489 -2326 3501
rect -2210 3898 -1948 3910
rect -2210 3501 -2204 3898
rect -1954 3501 -1948 3898
rect -2210 3489 -1948 3501
rect -1832 3898 -1570 3910
rect -1832 3501 -1826 3898
rect -1576 3501 -1570 3898
rect -1832 3489 -1570 3501
rect -1454 3898 -1192 3910
rect -1454 3501 -1448 3898
rect -1198 3501 -1192 3898
rect -1454 3489 -1192 3501
rect -1076 3898 -814 3910
rect -1076 3501 -1070 3898
rect -820 3501 -814 3898
rect -1076 3489 -814 3501
rect -698 3898 -436 3910
rect -698 3501 -692 3898
rect -442 3501 -436 3898
rect -698 3489 -436 3501
rect -320 3898 -58 3910
rect -320 3501 -314 3898
rect -64 3501 -58 3898
rect -320 3489 -58 3501
rect 58 3898 320 3910
rect 58 3501 64 3898
rect 314 3501 320 3898
rect 58 3489 320 3501
rect 436 3898 698 3910
rect 436 3501 442 3898
rect 692 3501 698 3898
rect 436 3489 698 3501
rect 814 3898 1076 3910
rect 814 3501 820 3898
rect 1070 3501 1076 3898
rect 814 3489 1076 3501
rect 1192 3898 1454 3910
rect 1192 3501 1198 3898
rect 1448 3501 1454 3898
rect 1192 3489 1454 3501
rect 1570 3898 1832 3910
rect 1570 3501 1576 3898
rect 1826 3501 1832 3898
rect 1570 3489 1832 3501
rect 1948 3898 2210 3910
rect 1948 3501 1954 3898
rect 2204 3501 2210 3898
rect 1948 3489 2210 3501
rect 2326 3898 2588 3910
rect 2326 3501 2332 3898
rect 2582 3501 2588 3898
rect 2326 3489 2588 3501
rect 2704 3898 2966 3910
rect 2704 3501 2710 3898
rect 2960 3501 2966 3898
rect 2704 3489 2966 3501
rect 3082 3898 3344 3910
rect 3082 3501 3088 3898
rect 3338 3501 3344 3898
rect 3082 3489 3344 3501
rect 3460 3898 3722 3910
rect 3460 3501 3466 3898
rect 3716 3501 3722 3898
rect 3460 3489 3722 3501
rect 3838 3898 4100 3910
rect 3838 3501 3844 3898
rect 4094 3501 4100 3898
rect 3838 3489 4100 3501
rect 4216 3898 4478 3910
rect 4216 3501 4222 3898
rect 4472 3501 4478 3898
rect 4216 3489 4478 3501
rect 4594 3898 4856 3910
rect 4594 3501 4600 3898
rect 4850 3501 4856 3898
rect 4594 3489 4856 3501
rect 4972 3898 5234 3910
rect 4972 3501 4978 3898
rect 5228 3501 5234 3898
rect 4972 3489 5234 3501
rect 5350 3898 5612 3910
rect 5350 3501 5356 3898
rect 5606 3501 5612 3898
rect 5350 3489 5612 3501
rect 5728 3898 5990 3910
rect 5728 3501 5734 3898
rect 5984 3501 5990 3898
rect 5728 3489 5990 3501
rect 6106 3898 6368 3910
rect 6106 3501 6112 3898
rect 6362 3501 6368 3898
rect 6106 3489 6368 3501
rect 6484 3898 6746 3910
rect 6484 3501 6490 3898
rect 6740 3501 6746 3898
rect 6484 3489 6746 3501
rect 6862 3898 7124 3910
rect 6862 3501 6868 3898
rect 7118 3501 7124 3898
rect 6862 3489 7124 3501
rect 7240 3898 7502 3910
rect 7240 3501 7246 3898
rect 7496 3501 7502 3898
rect 7240 3489 7502 3501
rect 7618 3898 7880 3910
rect 7618 3501 7624 3898
rect 7874 3501 7880 3898
rect 7618 3489 7880 3501
rect 7996 3898 8258 3910
rect 7996 3501 8002 3898
rect 8252 3501 8258 3898
rect 7996 3489 8258 3501
rect 8374 3898 8636 3910
rect 8374 3501 8380 3898
rect 8630 3501 8636 3898
rect 8374 3489 8636 3501
rect 8752 3898 9014 3910
rect 8752 3501 8758 3898
rect 9008 3501 9014 3898
rect 8752 3489 9014 3501
rect 9130 3898 9392 3910
rect 9130 3501 9136 3898
rect 9386 3501 9392 3898
rect 9130 3489 9392 3501
rect 9508 3898 9770 3910
rect 9508 3501 9514 3898
rect 9764 3501 9770 3898
rect 9508 3489 9770 3501
rect 9886 3898 10148 3910
rect 9886 3501 9892 3898
rect 10142 3501 10148 3898
rect 9886 3489 10148 3501
rect 10264 3898 10526 3910
rect 10264 3501 10270 3898
rect 10520 3501 10526 3898
rect 10264 3489 10526 3501
rect 10642 3898 10904 3910
rect 10642 3501 10648 3898
rect 10898 3501 10904 3898
rect 10642 3489 10904 3501
rect 11020 3898 11282 3910
rect 11020 3501 11026 3898
rect 11276 3501 11282 3898
rect 11020 3489 11282 3501
rect 11398 3898 11660 3910
rect 11398 3501 11404 3898
rect 11654 3501 11660 3898
rect 11398 3489 11660 3501
rect 11776 3898 12038 3910
rect 11776 3501 11782 3898
rect 12032 3501 12038 3898
rect 11776 3489 12038 3501
rect 12154 3898 12416 3910
rect 12154 3501 12160 3898
rect 12410 3501 12416 3898
rect 12154 3489 12416 3501
rect 12532 3898 12794 3910
rect 12532 3501 12538 3898
rect 12788 3501 12794 3898
rect 12532 3489 12794 3501
rect 12910 3898 13172 3910
rect 12910 3501 12916 3898
rect 13166 3501 13172 3898
rect 12910 3489 13172 3501
rect -13172 -3501 -12910 -3489
rect -13172 -3898 -13166 -3501
rect -12916 -3898 -12910 -3501
rect -13172 -3910 -12910 -3898
rect -12794 -3501 -12532 -3489
rect -12794 -3898 -12788 -3501
rect -12538 -3898 -12532 -3501
rect -12794 -3910 -12532 -3898
rect -12416 -3501 -12154 -3489
rect -12416 -3898 -12410 -3501
rect -12160 -3898 -12154 -3501
rect -12416 -3910 -12154 -3898
rect -12038 -3501 -11776 -3489
rect -12038 -3898 -12032 -3501
rect -11782 -3898 -11776 -3501
rect -12038 -3910 -11776 -3898
rect -11660 -3501 -11398 -3489
rect -11660 -3898 -11654 -3501
rect -11404 -3898 -11398 -3501
rect -11660 -3910 -11398 -3898
rect -11282 -3501 -11020 -3489
rect -11282 -3898 -11276 -3501
rect -11026 -3898 -11020 -3501
rect -11282 -3910 -11020 -3898
rect -10904 -3501 -10642 -3489
rect -10904 -3898 -10898 -3501
rect -10648 -3898 -10642 -3501
rect -10904 -3910 -10642 -3898
rect -10526 -3501 -10264 -3489
rect -10526 -3898 -10520 -3501
rect -10270 -3898 -10264 -3501
rect -10526 -3910 -10264 -3898
rect -10148 -3501 -9886 -3489
rect -10148 -3898 -10142 -3501
rect -9892 -3898 -9886 -3501
rect -10148 -3910 -9886 -3898
rect -9770 -3501 -9508 -3489
rect -9770 -3898 -9764 -3501
rect -9514 -3898 -9508 -3501
rect -9770 -3910 -9508 -3898
rect -9392 -3501 -9130 -3489
rect -9392 -3898 -9386 -3501
rect -9136 -3898 -9130 -3501
rect -9392 -3910 -9130 -3898
rect -9014 -3501 -8752 -3489
rect -9014 -3898 -9008 -3501
rect -8758 -3898 -8752 -3501
rect -9014 -3910 -8752 -3898
rect -8636 -3501 -8374 -3489
rect -8636 -3898 -8630 -3501
rect -8380 -3898 -8374 -3501
rect -8636 -3910 -8374 -3898
rect -8258 -3501 -7996 -3489
rect -8258 -3898 -8252 -3501
rect -8002 -3898 -7996 -3501
rect -8258 -3910 -7996 -3898
rect -7880 -3501 -7618 -3489
rect -7880 -3898 -7874 -3501
rect -7624 -3898 -7618 -3501
rect -7880 -3910 -7618 -3898
rect -7502 -3501 -7240 -3489
rect -7502 -3898 -7496 -3501
rect -7246 -3898 -7240 -3501
rect -7502 -3910 -7240 -3898
rect -7124 -3501 -6862 -3489
rect -7124 -3898 -7118 -3501
rect -6868 -3898 -6862 -3501
rect -7124 -3910 -6862 -3898
rect -6746 -3501 -6484 -3489
rect -6746 -3898 -6740 -3501
rect -6490 -3898 -6484 -3501
rect -6746 -3910 -6484 -3898
rect -6368 -3501 -6106 -3489
rect -6368 -3898 -6362 -3501
rect -6112 -3898 -6106 -3501
rect -6368 -3910 -6106 -3898
rect -5990 -3501 -5728 -3489
rect -5990 -3898 -5984 -3501
rect -5734 -3898 -5728 -3501
rect -5990 -3910 -5728 -3898
rect -5612 -3501 -5350 -3489
rect -5612 -3898 -5606 -3501
rect -5356 -3898 -5350 -3501
rect -5612 -3910 -5350 -3898
rect -5234 -3501 -4972 -3489
rect -5234 -3898 -5228 -3501
rect -4978 -3898 -4972 -3501
rect -5234 -3910 -4972 -3898
rect -4856 -3501 -4594 -3489
rect -4856 -3898 -4850 -3501
rect -4600 -3898 -4594 -3501
rect -4856 -3910 -4594 -3898
rect -4478 -3501 -4216 -3489
rect -4478 -3898 -4472 -3501
rect -4222 -3898 -4216 -3501
rect -4478 -3910 -4216 -3898
rect -4100 -3501 -3838 -3489
rect -4100 -3898 -4094 -3501
rect -3844 -3898 -3838 -3501
rect -4100 -3910 -3838 -3898
rect -3722 -3501 -3460 -3489
rect -3722 -3898 -3716 -3501
rect -3466 -3898 -3460 -3501
rect -3722 -3910 -3460 -3898
rect -3344 -3501 -3082 -3489
rect -3344 -3898 -3338 -3501
rect -3088 -3898 -3082 -3501
rect -3344 -3910 -3082 -3898
rect -2966 -3501 -2704 -3489
rect -2966 -3898 -2960 -3501
rect -2710 -3898 -2704 -3501
rect -2966 -3910 -2704 -3898
rect -2588 -3501 -2326 -3489
rect -2588 -3898 -2582 -3501
rect -2332 -3898 -2326 -3501
rect -2588 -3910 -2326 -3898
rect -2210 -3501 -1948 -3489
rect -2210 -3898 -2204 -3501
rect -1954 -3898 -1948 -3501
rect -2210 -3910 -1948 -3898
rect -1832 -3501 -1570 -3489
rect -1832 -3898 -1826 -3501
rect -1576 -3898 -1570 -3501
rect -1832 -3910 -1570 -3898
rect -1454 -3501 -1192 -3489
rect -1454 -3898 -1448 -3501
rect -1198 -3898 -1192 -3501
rect -1454 -3910 -1192 -3898
rect -1076 -3501 -814 -3489
rect -1076 -3898 -1070 -3501
rect -820 -3898 -814 -3501
rect -1076 -3910 -814 -3898
rect -698 -3501 -436 -3489
rect -698 -3898 -692 -3501
rect -442 -3898 -436 -3501
rect -698 -3910 -436 -3898
rect -320 -3501 -58 -3489
rect -320 -3898 -314 -3501
rect -64 -3898 -58 -3501
rect -320 -3910 -58 -3898
rect 58 -3501 320 -3489
rect 58 -3898 64 -3501
rect 314 -3898 320 -3501
rect 58 -3910 320 -3898
rect 436 -3501 698 -3489
rect 436 -3898 442 -3501
rect 692 -3898 698 -3501
rect 436 -3910 698 -3898
rect 814 -3501 1076 -3489
rect 814 -3898 820 -3501
rect 1070 -3898 1076 -3501
rect 814 -3910 1076 -3898
rect 1192 -3501 1454 -3489
rect 1192 -3898 1198 -3501
rect 1448 -3898 1454 -3501
rect 1192 -3910 1454 -3898
rect 1570 -3501 1832 -3489
rect 1570 -3898 1576 -3501
rect 1826 -3898 1832 -3501
rect 1570 -3910 1832 -3898
rect 1948 -3501 2210 -3489
rect 1948 -3898 1954 -3501
rect 2204 -3898 2210 -3501
rect 1948 -3910 2210 -3898
rect 2326 -3501 2588 -3489
rect 2326 -3898 2332 -3501
rect 2582 -3898 2588 -3501
rect 2326 -3910 2588 -3898
rect 2704 -3501 2966 -3489
rect 2704 -3898 2710 -3501
rect 2960 -3898 2966 -3501
rect 2704 -3910 2966 -3898
rect 3082 -3501 3344 -3489
rect 3082 -3898 3088 -3501
rect 3338 -3898 3344 -3501
rect 3082 -3910 3344 -3898
rect 3460 -3501 3722 -3489
rect 3460 -3898 3466 -3501
rect 3716 -3898 3722 -3501
rect 3460 -3910 3722 -3898
rect 3838 -3501 4100 -3489
rect 3838 -3898 3844 -3501
rect 4094 -3898 4100 -3501
rect 3838 -3910 4100 -3898
rect 4216 -3501 4478 -3489
rect 4216 -3898 4222 -3501
rect 4472 -3898 4478 -3501
rect 4216 -3910 4478 -3898
rect 4594 -3501 4856 -3489
rect 4594 -3898 4600 -3501
rect 4850 -3898 4856 -3501
rect 4594 -3910 4856 -3898
rect 4972 -3501 5234 -3489
rect 4972 -3898 4978 -3501
rect 5228 -3898 5234 -3501
rect 4972 -3910 5234 -3898
rect 5350 -3501 5612 -3489
rect 5350 -3898 5356 -3501
rect 5606 -3898 5612 -3501
rect 5350 -3910 5612 -3898
rect 5728 -3501 5990 -3489
rect 5728 -3898 5734 -3501
rect 5984 -3898 5990 -3501
rect 5728 -3910 5990 -3898
rect 6106 -3501 6368 -3489
rect 6106 -3898 6112 -3501
rect 6362 -3898 6368 -3501
rect 6106 -3910 6368 -3898
rect 6484 -3501 6746 -3489
rect 6484 -3898 6490 -3501
rect 6740 -3898 6746 -3501
rect 6484 -3910 6746 -3898
rect 6862 -3501 7124 -3489
rect 6862 -3898 6868 -3501
rect 7118 -3898 7124 -3501
rect 6862 -3910 7124 -3898
rect 7240 -3501 7502 -3489
rect 7240 -3898 7246 -3501
rect 7496 -3898 7502 -3501
rect 7240 -3910 7502 -3898
rect 7618 -3501 7880 -3489
rect 7618 -3898 7624 -3501
rect 7874 -3898 7880 -3501
rect 7618 -3910 7880 -3898
rect 7996 -3501 8258 -3489
rect 7996 -3898 8002 -3501
rect 8252 -3898 8258 -3501
rect 7996 -3910 8258 -3898
rect 8374 -3501 8636 -3489
rect 8374 -3898 8380 -3501
rect 8630 -3898 8636 -3501
rect 8374 -3910 8636 -3898
rect 8752 -3501 9014 -3489
rect 8752 -3898 8758 -3501
rect 9008 -3898 9014 -3501
rect 8752 -3910 9014 -3898
rect 9130 -3501 9392 -3489
rect 9130 -3898 9136 -3501
rect 9386 -3898 9392 -3501
rect 9130 -3910 9392 -3898
rect 9508 -3501 9770 -3489
rect 9508 -3898 9514 -3501
rect 9764 -3898 9770 -3501
rect 9508 -3910 9770 -3898
rect 9886 -3501 10148 -3489
rect 9886 -3898 9892 -3501
rect 10142 -3898 10148 -3501
rect 9886 -3910 10148 -3898
rect 10264 -3501 10526 -3489
rect 10264 -3898 10270 -3501
rect 10520 -3898 10526 -3501
rect 10264 -3910 10526 -3898
rect 10642 -3501 10904 -3489
rect 10642 -3898 10648 -3501
rect 10898 -3898 10904 -3501
rect 10642 -3910 10904 -3898
rect 11020 -3501 11282 -3489
rect 11020 -3898 11026 -3501
rect 11276 -3898 11282 -3501
rect 11020 -3910 11282 -3898
rect 11398 -3501 11660 -3489
rect 11398 -3898 11404 -3501
rect 11654 -3898 11660 -3501
rect 11398 -3910 11660 -3898
rect 11776 -3501 12038 -3489
rect 11776 -3898 11782 -3501
rect 12032 -3898 12038 -3501
rect 11776 -3910 12038 -3898
rect 12154 -3501 12416 -3489
rect 12154 -3898 12160 -3501
rect 12410 -3898 12416 -3501
rect 12154 -3910 12416 -3898
rect 12532 -3501 12794 -3489
rect 12532 -3898 12538 -3501
rect 12788 -3898 12794 -3501
rect 12532 -3910 12794 -3898
rect 12910 -3501 13172 -3489
rect 12910 -3898 12916 -3501
rect 13166 -3898 13172 -3501
rect 12910 -3910 13172 -3898
<< properties >>
string FIXED_BBOX -13295 -4029 13295 4029
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 35 m 1 nx 70 wmin 1.410 lmin 0.50 rho 2000 val 49.912k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

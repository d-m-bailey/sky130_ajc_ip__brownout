magic
tech sky130A
magscale 1 2
timestamp 1712463840
<< metal4 >>
rect -3349 19039 3349 19080
rect -3349 12961 3093 19039
rect 3329 12961 3349 19039
rect -3349 12920 3349 12961
rect -3349 12639 3349 12680
rect -3349 6561 3093 12639
rect 3329 6561 3349 12639
rect -3349 6520 3349 6561
rect -3349 6239 3349 6280
rect -3349 161 3093 6239
rect 3329 161 3349 6239
rect -3349 120 3349 161
rect -3349 -161 3349 -120
rect -3349 -6239 3093 -161
rect 3329 -6239 3349 -161
rect -3349 -6280 3349 -6239
rect -3349 -6561 3349 -6520
rect -3349 -12639 3093 -6561
rect 3329 -12639 3349 -6561
rect -3349 -12680 3349 -12639
rect -3349 -12961 3349 -12920
rect -3349 -19039 3093 -12961
rect 3329 -19039 3349 -12961
rect -3349 -19080 3349 -19039
<< via4 >>
rect 3093 12961 3329 19039
rect 3093 6561 3329 12639
rect 3093 161 3329 6239
rect 3093 -6239 3329 -161
rect 3093 -12639 3329 -6561
rect 3093 -19039 3329 -12961
<< mimcap2 >>
rect -3269 18960 2731 19000
rect -3269 13040 -3229 18960
rect 2691 13040 2731 18960
rect -3269 13000 2731 13040
rect -3269 12560 2731 12600
rect -3269 6640 -3229 12560
rect 2691 6640 2731 12560
rect -3269 6600 2731 6640
rect -3269 6160 2731 6200
rect -3269 240 -3229 6160
rect 2691 240 2731 6160
rect -3269 200 2731 240
rect -3269 -240 2731 -200
rect -3269 -6160 -3229 -240
rect 2691 -6160 2731 -240
rect -3269 -6200 2731 -6160
rect -3269 -6640 2731 -6600
rect -3269 -12560 -3229 -6640
rect 2691 -12560 2731 -6640
rect -3269 -12600 2731 -12560
rect -3269 -13040 2731 -13000
rect -3269 -18960 -3229 -13040
rect 2691 -18960 2731 -13040
rect -3269 -19000 2731 -18960
<< mimcap2contact >>
rect -3229 13040 2691 18960
rect -3229 6640 2691 12560
rect -3229 240 2691 6160
rect -3229 -6160 2691 -240
rect -3229 -12560 2691 -6640
rect -3229 -18960 2691 -13040
<< metal5 >>
rect -429 18984 -109 19200
rect 3051 19039 3371 19200
rect -3253 18960 2715 18984
rect -3253 13040 -3229 18960
rect 2691 13040 2715 18960
rect -3253 13016 2715 13040
rect -429 12584 -109 13016
rect 3051 12961 3093 19039
rect 3329 12961 3371 19039
rect 3051 12639 3371 12961
rect -3253 12560 2715 12584
rect -3253 6640 -3229 12560
rect 2691 6640 2715 12560
rect -3253 6616 2715 6640
rect -429 6184 -109 6616
rect 3051 6561 3093 12639
rect 3329 6561 3371 12639
rect 3051 6239 3371 6561
rect -3253 6160 2715 6184
rect -3253 240 -3229 6160
rect 2691 240 2715 6160
rect -3253 216 2715 240
rect -429 -216 -109 216
rect 3051 161 3093 6239
rect 3329 161 3371 6239
rect 3051 -161 3371 161
rect -3253 -240 2715 -216
rect -3253 -6160 -3229 -240
rect 2691 -6160 2715 -240
rect -3253 -6184 2715 -6160
rect -429 -6616 -109 -6184
rect 3051 -6239 3093 -161
rect 3329 -6239 3371 -161
rect 3051 -6561 3371 -6239
rect -3253 -6640 2715 -6616
rect -3253 -12560 -3229 -6640
rect 2691 -12560 2715 -6640
rect -3253 -12584 2715 -12560
rect -429 -13016 -109 -12584
rect 3051 -12639 3093 -6561
rect 3329 -12639 3371 -6561
rect 3051 -12961 3371 -12639
rect -3253 -13040 2715 -13016
rect -3253 -18960 -3229 -13040
rect 2691 -18960 2715 -13040
rect -3253 -18984 2715 -18960
rect -429 -19200 -109 -18984
rect 3051 -19039 3093 -12961
rect 3329 -19039 3371 -12961
rect 3051 -19200 3371 -19039
<< properties >>
string FIXED_BBOX -3349 12920 2811 19080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

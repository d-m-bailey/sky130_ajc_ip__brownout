magic
tech sky130A
magscale 1 2
timestamp 1712709231
<< pwell >>
rect -307 -25050 307 25050
<< psubdiff >>
rect -271 24980 -175 25014
rect 175 24980 271 25014
rect -271 24918 -237 24980
rect 237 24918 271 24980
rect -271 -24980 -237 -24918
rect 237 -24980 271 -24918
rect -271 -25014 -175 -24980
rect 175 -25014 271 -24980
<< psubdiffcont >>
rect -175 24980 175 25014
rect -271 -24918 -237 24918
rect 237 -24918 271 24918
rect -175 -25014 175 -24980
<< xpolycontact >>
rect -141 24452 141 24884
rect -141 52 141 484
rect -141 -484 141 -52
rect -141 -24884 141 -24452
<< xpolyres >>
rect -141 484 141 24452
rect -141 -24452 141 -484
<< locali >>
rect -271 24980 -175 25014
rect 175 24980 271 25014
rect -271 24918 -237 24980
rect 237 24918 271 24980
rect -271 -24980 -237 -24918
rect 237 -24980 271 -24918
rect -271 -25014 -175 -24980
rect 175 -25014 271 -24980
<< viali >>
rect -125 24469 125 24866
rect -125 70 125 467
rect -125 -467 125 -70
rect -125 -24866 125 -24469
<< metal1 >>
rect -131 24866 131 24878
rect -131 24469 -125 24866
rect 125 24469 131 24866
rect -131 24457 131 24469
rect -131 467 131 479
rect -131 70 -125 467
rect 125 70 131 467
rect -131 58 131 70
rect -131 -70 131 -58
rect -131 -467 -125 -70
rect 125 -467 131 -70
rect -131 -479 131 -467
rect -131 -24469 131 -24457
rect -131 -24866 -125 -24469
rect 125 -24866 131 -24469
rect -131 -24878 131 -24866
<< properties >>
string FIXED_BBOX -254 -24997 254 24997
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 120 m 2 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 170.479k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

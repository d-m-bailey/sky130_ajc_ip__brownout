magic
tech sky130A
magscale 1 2
timestamp 1712901446
<< error_s >>
rect 39827 23173 39828 23227
rect 39887 23123 39888 23173
rect 39887 22853 39888 22937
<< pwell >>
rect -1182 40391 42901 40527
rect -1182 -559 -1046 40391
rect 42765 -559 42901 40391
rect -1182 -695 42901 -559
<< psubdiff >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< psubdiffcont >>
rect -1086 40457 42805 40491
rect -1146 -599 -1112 40431
rect 42831 -599 42865 40431
rect -1086 -659 42805 -625
<< locali >>
rect 41825 62329 41873 62377
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< viali >>
rect -1086 40457 42805 40491
rect -1146 -556 -1112 40404
rect 42831 -567 42865 40393
rect -1086 -659 42805 -625
<< metal1 >>
rect -1186 40491 42905 40531
rect -1186 40457 -1086 40491
rect 42805 40457 42905 40491
rect -1186 40404 42905 40457
rect -1186 -556 -1146 40404
rect -1112 40393 42905 40404
rect -1112 40391 42831 40393
rect -1112 -556 -1046 40391
rect -1186 -559 -1046 -556
rect 42765 -559 42831 40391
rect -1186 -567 42831 -559
rect 42865 -567 42905 40393
rect -1186 -625 42905 -567
rect -1186 -659 -1086 -625
rect 42805 -659 42905 -625
rect -1186 -699 42905 -659
<< metal2 >>
rect 31111 38144 31167 38151
rect 38119 38144 38197 38153
rect 31109 38142 31169 38144
rect 31109 38086 31111 38142
rect 31167 38086 31169 38142
rect 30945 37995 31001 38002
rect 30943 37993 31003 37995
rect 30943 37937 30945 37993
rect 31001 37937 31003 37993
rect 30810 37852 30866 37859
rect 30808 37850 30868 37852
rect 30808 37794 30810 37850
rect 30866 37794 30868 37850
rect 30657 37703 30713 37710
rect 30655 37701 30715 37703
rect 30655 37645 30657 37701
rect 30713 37645 30715 37701
rect 30112 37569 30168 37576
rect 30110 37567 30170 37569
rect 30110 37511 30112 37567
rect 30168 37511 30170 37567
rect 29963 35081 30019 35088
rect 29961 35079 30021 35081
rect 29961 35023 29963 35079
rect 30019 35023 30021 35079
rect 19684 34398 19744 34407
rect 15261 4203 15317 4210
rect 15259 4201 15319 4203
rect 15259 4145 15261 4201
rect 15317 4145 15319 4201
rect 15259 3495 15319 4145
rect 15157 3435 15319 3495
rect 18496 3531 18556 3540
rect 19684 3529 19744 34338
rect 24320 30877 24380 30886
rect 19930 28201 19990 28210
rect 19921 28141 19930 28197
rect 19990 28141 19999 28197
rect 19930 4203 19990 28141
rect 21332 27822 21388 27829
rect 21330 27820 21390 27822
rect 21330 27764 21332 27820
rect 21388 27764 21390 27820
rect 21330 23716 21390 27764
rect 23126 27660 23182 27667
rect 23124 27658 23184 27660
rect 23124 27602 23126 27658
rect 23182 27602 23184 27658
rect 21508 26814 21564 26821
rect 21506 26812 21566 26814
rect 21506 26756 21508 26812
rect 21564 26756 21566 26812
rect 21506 22328 21566 26756
rect 23124 23396 23184 27602
rect 23637 26947 23693 26954
rect 23635 26945 23695 26947
rect 23635 26889 23637 26945
rect 23693 26889 23695 26945
rect 23635 23875 23695 26889
rect 24320 26680 24380 30817
rect 29742 30313 29802 30322
rect 26802 30024 26858 30033
rect 26802 29959 26858 29968
rect 27842 30026 27902 30035
rect 26785 28398 26845 28407
rect 26785 28329 26845 28338
rect 26787 27893 26843 28329
rect 27842 28044 27902 29966
rect 29742 28396 29802 30253
rect 29742 28340 29744 28396
rect 29800 28340 29802 28396
rect 29742 28338 29802 28340
rect 29744 28331 29800 28338
rect 27842 27988 27844 28044
rect 27900 27988 27902 28044
rect 27842 27986 27902 27988
rect 27844 27979 27900 27986
rect 26787 27837 26932 27893
rect 25396 27508 25452 27515
rect 24320 26624 24322 26680
rect 24378 26624 24380 26680
rect 24320 26622 24380 26624
rect 25394 27506 25454 27508
rect 25394 27450 25396 27506
rect 25452 27450 25454 27506
rect 24322 26615 24378 26622
rect 23448 23815 23695 23875
rect 23124 23336 23498 23396
rect 21337 22268 21566 22328
rect 21337 22054 21397 22268
rect 23438 22074 23498 23336
rect 25394 22642 25454 27450
rect 27504 27368 27560 27375
rect 27502 27366 27562 27368
rect 27502 27310 27504 27366
rect 27560 27310 27562 27366
rect 25556 27228 25612 27235
rect 25554 27226 25614 27228
rect 25554 27170 25556 27226
rect 25612 27170 25614 27226
rect 25554 23786 25614 27170
rect 25394 22582 25614 22642
rect 25554 22032 25614 22582
rect 27502 22332 27562 27310
rect 27676 27088 27732 27095
rect 27674 27086 27734 27088
rect 27674 27030 27676 27086
rect 27732 27030 27734 27086
rect 27674 23750 27734 27030
rect 29961 25717 30021 35023
rect 29961 25648 30021 25657
rect 29783 23848 29839 23857
rect 29783 23783 29839 23792
rect 29776 22335 29832 22342
rect 30110 22335 30170 37511
rect 30502 37443 30558 37450
rect 30500 37441 30560 37443
rect 30500 37385 30502 37441
rect 30558 37385 30560 37441
rect 30266 37312 30322 37319
rect 30264 37310 30324 37312
rect 30264 37254 30266 37310
rect 30322 37254 30324 37310
rect 30264 23850 30324 37254
rect 30383 37187 30439 37194
rect 30264 23781 30324 23790
rect 30381 37185 30441 37187
rect 30381 37129 30383 37185
rect 30439 37129 30441 37185
rect 29774 22333 29834 22335
rect 27502 22272 27726 22332
rect 27666 22088 27726 22272
rect 29774 22277 29776 22333
rect 29832 22277 29834 22333
rect 29774 22108 29834 22277
rect 30110 22266 30170 22275
rect 30381 22306 30441 37129
rect 30500 26524 30560 37385
rect 30500 26455 30560 26464
rect 30655 26370 30715 37645
rect 30655 26301 30715 26310
rect 30808 26202 30868 37794
rect 30808 26133 30868 26142
rect 30943 26029 31003 37937
rect 30943 25960 31003 25969
rect 31109 25870 31169 38086
rect 38119 38084 38128 38144
rect 38188 38084 38197 38144
rect 38119 38075 38197 38084
rect 37475 37995 37553 38004
rect 37475 37935 37484 37995
rect 37544 37935 37553 37995
rect 37475 37926 37553 37935
rect 36831 37792 36840 37852
rect 36900 37792 36909 37852
rect 36187 37703 36265 37712
rect 36187 37643 36196 37703
rect 36256 37643 36265 37703
rect 36187 37634 36265 37643
rect 35543 37569 35621 37578
rect 35543 37509 35552 37569
rect 35612 37509 35621 37569
rect 35543 37500 35621 37509
rect 34908 37443 34968 37452
rect 34908 37374 34968 37383
rect 34255 37312 34333 37321
rect 34255 37252 34264 37312
rect 34324 37252 34333 37312
rect 34255 37243 34333 37252
rect 33611 37187 33689 37196
rect 33611 37127 33620 37187
rect 33680 37127 33689 37187
rect 33611 37118 33689 37127
rect 40462 33036 40536 33045
rect 40462 32980 40471 33036
rect 40527 32980 40536 33036
rect 40462 32975 40536 32980
rect 40469 32578 40529 32975
rect 40377 32518 40529 32578
rect 40377 32187 40437 32518
rect 40767 32358 40823 32365
rect 40765 32356 40825 32358
rect 40765 32300 40767 32356
rect 40823 32300 40825 32356
rect 40377 32127 40495 32187
rect 40293 30996 40367 31005
rect 40293 30940 40302 30996
rect 40358 30940 40367 30996
rect 40293 30935 40367 30940
rect 40300 28201 40360 30935
rect 40300 28132 40360 28141
rect 34908 27822 34968 27831
rect 34908 27753 34968 27762
rect 34255 27600 34264 27660
rect 34324 27600 34333 27660
rect 34924 27586 34952 27753
rect 37208 27508 37268 27517
rect 37208 27439 37268 27448
rect 37224 27368 37252 27439
rect 37484 27368 37544 27377
rect 37484 27299 37544 27308
rect 37500 27224 37528 27299
rect 38119 27168 38128 27228
rect 38188 27168 38197 27228
rect 38763 27088 38841 27097
rect 38763 27028 38772 27088
rect 38832 27028 38841 27088
rect 38763 27019 38841 27028
rect 39432 26956 39460 27250
rect 39416 26947 39476 26956
rect 39416 26878 39476 26887
rect 40076 26823 40104 27022
rect 40060 26814 40120 26823
rect 40060 26745 40120 26754
rect 40435 26682 40495 32127
rect 40765 28046 40825 32300
rect 40765 27977 40825 27986
rect 40435 26613 40495 26622
rect 33243 26524 33299 26531
rect 33241 26522 33301 26524
rect 33241 26466 33243 26522
rect 33299 26466 33301 26522
rect 31897 25870 31953 25877
rect 31109 25801 31169 25810
rect 31895 25868 31955 25870
rect 31895 25812 31897 25868
rect 31953 25812 31955 25868
rect 31895 23786 31955 25812
rect 33241 22898 33301 26466
rect 35943 26370 35999 26377
rect 35941 26368 36001 26370
rect 35941 26312 35943 26368
rect 35999 26312 36001 26368
rect 34007 26202 34063 26209
rect 34005 26200 34065 26202
rect 34005 26144 34007 26200
rect 34063 26144 34065 26200
rect 34005 23812 34065 26144
rect 33241 22838 33465 22898
rect 35941 22315 36001 26312
rect 36128 26027 36188 26029
rect 36121 25971 36130 26027
rect 36186 25971 36195 26027
rect 36128 23792 36188 25971
rect 38020 25717 38076 25724
rect 38018 25715 38078 25717
rect 38018 25659 38020 25715
rect 38076 25659 38078 25715
rect 31892 22306 31948 22313
rect 30381 22237 30441 22246
rect 31890 22304 31950 22306
rect 31890 22248 31892 22304
rect 31948 22248 31950 22304
rect 35941 22255 36175 22315
rect 31890 22097 31950 22248
rect 36115 22040 36175 22255
rect 38018 22281 38078 25659
rect 38018 22221 38276 22281
rect 38216 22103 38276 22221
rect 19930 4134 19990 4143
rect 19677 3473 19686 3529
rect 19742 3473 19751 3529
rect 19684 3471 19744 3473
rect 18496 3462 18556 3471
<< via2 >>
rect 31111 38086 31167 38142
rect 30945 37937 31001 37993
rect 30810 37794 30866 37850
rect 30657 37645 30713 37701
rect 30112 37511 30168 37567
rect 29963 35023 30019 35079
rect 19684 34338 19744 34398
rect 15261 4145 15317 4201
rect 18496 3471 18556 3531
rect 24320 30817 24380 30877
rect 19930 28141 19990 28201
rect 21332 27764 21388 27820
rect 23126 27602 23182 27658
rect 21508 26756 21564 26812
rect 23637 26889 23693 26945
rect 29742 30253 29802 30313
rect 26802 29968 26858 30024
rect 27842 29966 27902 30026
rect 26785 28338 26845 28398
rect 29744 28340 29800 28396
rect 27844 27988 27900 28044
rect 24322 26624 24378 26680
rect 25396 27450 25452 27506
rect 27504 27310 27560 27366
rect 25556 27170 25612 27226
rect 27676 27030 27732 27086
rect 29961 25657 30021 25717
rect 29783 23792 29839 23848
rect 30502 37385 30558 37441
rect 30266 37254 30322 37310
rect 30264 23790 30324 23850
rect 30383 37129 30439 37185
rect 29776 22277 29832 22333
rect 30110 22275 30170 22335
rect 30500 26464 30560 26524
rect 30655 26310 30715 26370
rect 30808 26142 30868 26202
rect 30943 25969 31003 26029
rect 38128 38084 38188 38144
rect 37484 37935 37544 37995
rect 36840 37792 36900 37852
rect 36196 37643 36256 37703
rect 35552 37509 35612 37569
rect 34908 37383 34968 37443
rect 34264 37252 34324 37312
rect 33620 37127 33680 37187
rect 40471 32980 40527 33036
rect 40767 32300 40823 32356
rect 40302 30940 40358 30996
rect 40300 28141 40360 28201
rect 34908 27762 34968 27822
rect 34264 27600 34324 27660
rect 37208 27448 37268 27508
rect 37484 27308 37544 27368
rect 38128 27168 38188 27228
rect 38772 27028 38832 27088
rect 39416 26887 39476 26947
rect 40060 26754 40120 26814
rect 40765 27986 40825 28046
rect 40435 26622 40495 26682
rect 33243 26466 33299 26522
rect 31109 25810 31169 25870
rect 31897 25812 31953 25868
rect 35943 26312 35999 26368
rect 34007 26144 34063 26200
rect 36130 25971 36186 26027
rect 38020 25659 38076 25715
rect 30381 22246 30441 22306
rect 31892 22248 31948 22304
rect 19930 4143 19990 4203
rect 19686 3473 19742 3529
<< metal3 >>
rect -44 75676 44853 75682
rect -44 75288 -38 75676
rect 350 75288 44459 75676
rect 44847 75288 44853 75676
rect -44 75282 44853 75288
rect -44 75216 44853 75222
rect -44 74828 422 75216
rect 810 74828 43999 75216
rect 44387 74828 44853 75216
rect -44 74822 44853 74828
rect -44 74756 44853 74762
rect -44 74368 882 74756
rect 1270 74368 43539 74756
rect 43927 74368 44853 74756
rect -44 74362 44853 74368
rect -44 74296 44853 74302
rect -44 73908 1342 74296
rect 1730 73908 43079 74296
rect 43467 73908 44853 74296
rect -44 73902 44853 73908
rect 2507 73892 2917 73902
rect -44 46187 44853 46193
rect -44 45799 1342 46187
rect 1730 45799 43079 46187
rect 43467 45799 44853 46187
rect -44 45793 44853 45799
rect -44 45727 44853 45733
rect -44 45339 882 45727
rect 1270 45339 43539 45727
rect 43927 45339 44853 45727
rect -44 45333 44853 45339
rect -44 45267 44853 45273
rect -44 44879 422 45267
rect 810 44879 43999 45267
rect 44387 44879 44853 45267
rect -44 44873 44853 44879
rect -44 44807 44853 44813
rect -44 44419 -38 44807
rect 350 44419 44459 44807
rect 44847 44419 44853 44807
rect -44 44413 44853 44419
rect 31106 38144 31172 38147
rect 38123 38144 38193 38149
rect 31106 38142 38128 38144
rect 31106 38086 31111 38142
rect 31167 38086 38128 38142
rect 31106 38084 38128 38086
rect 38188 38084 38193 38144
rect 31106 38081 31172 38084
rect 38123 38079 38193 38084
rect 30940 37995 31006 37998
rect 37479 37995 37549 38000
rect 30940 37993 37484 37995
rect 30940 37937 30945 37993
rect 31001 37937 37484 37993
rect 30940 37935 37484 37937
rect 37544 37935 37549 37995
rect 30940 37932 31006 37935
rect 37479 37930 37549 37935
rect 30805 37852 30871 37855
rect 36835 37852 36905 37857
rect 30805 37850 36840 37852
rect 30805 37794 30810 37850
rect 30866 37794 36840 37850
rect 30805 37792 36840 37794
rect 36900 37792 36905 37852
rect 30805 37789 30871 37792
rect 36835 37787 36905 37792
rect 30652 37703 30718 37706
rect 36191 37703 36261 37708
rect 30652 37701 36196 37703
rect 30652 37645 30657 37701
rect 30713 37645 36196 37701
rect 30652 37643 36196 37645
rect 36256 37643 36261 37703
rect 30652 37640 30718 37643
rect 36191 37638 36261 37643
rect 30107 37569 30173 37572
rect 35547 37569 35617 37574
rect 30107 37567 35552 37569
rect 30107 37511 30112 37567
rect 30168 37511 35552 37567
rect 30107 37509 35552 37511
rect 35612 37509 35617 37569
rect 30107 37506 30173 37509
rect 35547 37504 35617 37509
rect 30497 37443 30563 37446
rect 34903 37443 34973 37448
rect 30497 37441 34908 37443
rect 30497 37385 30502 37441
rect 30558 37385 34908 37441
rect 30497 37383 34908 37385
rect 34968 37383 34973 37443
rect 30497 37380 30563 37383
rect 34903 37378 34973 37383
rect 30261 37312 30327 37315
rect 34259 37312 34329 37317
rect 30261 37310 34264 37312
rect 30261 37254 30266 37310
rect 30322 37254 34264 37310
rect 30261 37252 34264 37254
rect 34324 37252 34329 37312
rect 30261 37249 30327 37252
rect 34259 37247 34329 37252
rect 30378 37187 30444 37190
rect 33615 37187 33685 37192
rect 30378 37185 33620 37187
rect 30378 37129 30383 37185
rect 30439 37129 33620 37185
rect 30378 37127 33620 37129
rect 33680 37127 33685 37187
rect 30378 37124 30444 37127
rect 33615 37122 33685 37127
rect 29958 35081 30024 35084
rect 29958 35079 30384 35081
rect 29958 35023 29963 35079
rect 30019 35075 30384 35079
rect 30019 35023 31282 35075
rect 29958 35021 31282 35023
rect 29958 35018 30024 35021
rect 19679 34398 19749 34403
rect 19679 34338 19684 34398
rect 19744 34338 30674 34398
rect 19679 34333 19749 34338
rect 40466 33036 40532 33041
rect 40466 32980 40471 33036
rect 40527 32980 40532 33036
rect 40466 32975 40532 32980
rect 40762 32358 40828 32361
rect 40633 32356 40828 32358
rect 40633 32300 40767 32356
rect 40823 32300 40828 32356
rect 40633 32298 40828 32300
rect 40762 32295 40828 32298
rect 40297 30996 40363 31001
rect 40297 30940 40302 30996
rect 40358 30940 40363 30996
rect 40297 30935 40363 30940
rect 24315 30877 24385 30882
rect 24315 30817 24320 30877
rect 24380 30817 25001 30877
rect 24315 30812 24385 30817
rect 29737 30313 29807 30318
rect 29737 30253 29742 30313
rect 29802 30253 30759 30313
rect 29737 30248 29807 30253
rect 26797 30026 26863 30029
rect 27837 30026 27907 30031
rect 26797 30024 27842 30026
rect 26797 29968 26802 30024
rect 26858 29968 27842 30024
rect 26797 29966 27842 29968
rect 27902 29966 27907 30026
rect 26797 29963 26863 29966
rect 27837 29961 27907 29966
rect 26780 28398 26850 28403
rect 29739 28398 29805 28401
rect 26780 28338 26785 28398
rect 26845 28396 29805 28398
rect 26845 28340 29744 28396
rect 29800 28340 29805 28396
rect 26845 28338 29805 28340
rect 26780 28333 26850 28338
rect 29739 28335 29805 28338
rect 19925 28201 19995 28206
rect 40295 28201 40365 28206
rect 19925 28141 19930 28201
rect 19990 28141 40300 28201
rect 40360 28141 40365 28201
rect 19925 28136 19995 28141
rect 40295 28136 40365 28141
rect 27839 28046 27905 28049
rect 40760 28046 40830 28051
rect 27839 28044 40765 28046
rect 27839 27988 27844 28044
rect 27900 27988 40765 28044
rect 27839 27986 40765 27988
rect 40825 27986 40830 28046
rect 27839 27983 27905 27986
rect 40760 27981 40830 27986
rect 21327 27822 21393 27825
rect 34903 27822 34973 27827
rect 21327 27820 34908 27822
rect 21327 27764 21332 27820
rect 21388 27764 34908 27820
rect 21327 27762 34908 27764
rect 34968 27762 34973 27822
rect 21327 27759 21393 27762
rect 34903 27757 34973 27762
rect 23121 27660 23187 27663
rect 34259 27660 34329 27665
rect 23121 27658 34264 27660
rect 23121 27602 23126 27658
rect 23182 27602 34264 27658
rect 23121 27600 34264 27602
rect 34324 27600 34329 27660
rect 23121 27597 23187 27600
rect 34259 27595 34329 27600
rect 25391 27508 25457 27511
rect 37203 27508 37273 27513
rect 25391 27506 37208 27508
rect 25391 27450 25396 27506
rect 25452 27450 37208 27506
rect 25391 27448 37208 27450
rect 37268 27448 37273 27508
rect 25391 27445 25457 27448
rect 37203 27443 37273 27448
rect 27499 27368 27565 27371
rect 37479 27368 37549 27373
rect 27499 27366 37484 27368
rect 27499 27310 27504 27366
rect 27560 27310 37484 27366
rect 27499 27308 37484 27310
rect 37544 27308 37549 27368
rect 27499 27305 27565 27308
rect 37479 27303 37549 27308
rect 25551 27228 25617 27231
rect 38123 27228 38193 27233
rect 25551 27226 38128 27228
rect 25551 27170 25556 27226
rect 25612 27170 38128 27226
rect 25551 27168 38128 27170
rect 38188 27168 38193 27228
rect 25551 27165 25617 27168
rect 38123 27163 38193 27168
rect 27671 27088 27737 27091
rect 38767 27088 38837 27093
rect 27671 27086 38772 27088
rect 27671 27030 27676 27086
rect 27732 27030 38772 27086
rect 27671 27028 38772 27030
rect 38832 27028 38837 27088
rect 27671 27025 27737 27028
rect 38767 27023 38837 27028
rect 23632 26947 23698 26950
rect 39411 26947 39481 26952
rect 23632 26945 39416 26947
rect 23632 26889 23637 26945
rect 23693 26889 39416 26945
rect 23632 26887 39416 26889
rect 39476 26887 39481 26947
rect 23632 26884 23698 26887
rect 39411 26882 39481 26887
rect 21503 26814 21569 26817
rect 40055 26814 40125 26819
rect 21503 26812 40060 26814
rect 21503 26756 21508 26812
rect 21564 26756 40060 26812
rect 21503 26754 40060 26756
rect 40120 26754 40125 26814
rect 21503 26751 21569 26754
rect 40055 26749 40125 26754
rect 24317 26682 24383 26685
rect 40430 26682 40500 26687
rect 24317 26680 40435 26682
rect 24317 26624 24322 26680
rect 24378 26624 40435 26680
rect 24317 26622 40435 26624
rect 40495 26622 40500 26682
rect 24317 26619 24383 26622
rect 40430 26617 40500 26622
rect 30495 26524 30565 26529
rect 33238 26524 33304 26527
rect 30495 26464 30500 26524
rect 30560 26522 33304 26524
rect 30560 26466 33243 26522
rect 33299 26466 33304 26522
rect 30560 26464 33304 26466
rect 30495 26459 30565 26464
rect 33238 26461 33304 26464
rect 30650 26370 30720 26375
rect 35938 26370 36004 26373
rect 30650 26310 30655 26370
rect 30715 26368 36004 26370
rect 30715 26312 35943 26368
rect 35999 26312 36004 26368
rect 30715 26310 36004 26312
rect 30650 26305 30720 26310
rect 35938 26307 36004 26310
rect 30803 26202 30873 26207
rect 34002 26202 34068 26205
rect 30803 26142 30808 26202
rect 30868 26200 34068 26202
rect 30868 26144 34007 26200
rect 34063 26144 34068 26200
rect 30868 26142 34068 26144
rect 30803 26137 30873 26142
rect 34002 26139 34068 26142
rect 30938 26029 31008 26034
rect 36125 26029 36191 26032
rect 30938 25969 30943 26029
rect 31003 26027 36191 26029
rect 31003 25971 36130 26027
rect 36186 25971 36191 26027
rect 31003 25969 36191 25971
rect 30938 25964 31008 25969
rect 36125 25966 36191 25969
rect 31104 25870 31174 25875
rect 31892 25870 31958 25873
rect 31104 25810 31109 25870
rect 31169 25868 31958 25870
rect 31169 25812 31897 25868
rect 31953 25812 31958 25868
rect 31169 25810 31958 25812
rect 31104 25805 31174 25810
rect 31892 25807 31958 25810
rect 29956 25717 30026 25722
rect 38015 25717 38081 25720
rect 29956 25657 29961 25717
rect 30021 25715 38081 25717
rect 30021 25659 38020 25715
rect 38076 25659 38081 25715
rect 30021 25657 38081 25659
rect 29956 25652 30026 25657
rect 38015 25654 38081 25657
rect 29778 23850 29844 23853
rect 30259 23850 30329 23855
rect 29778 23848 30264 23850
rect 29778 23792 29783 23848
rect 29839 23792 30264 23848
rect 29778 23790 30264 23792
rect 30324 23790 30329 23850
rect 29778 23787 29844 23790
rect 30259 23785 30329 23790
rect 29771 22335 29837 22338
rect 30105 22335 30175 22340
rect 29771 22333 30110 22335
rect 29771 22277 29776 22333
rect 29832 22277 30110 22333
rect 29771 22275 30110 22277
rect 30170 22275 30175 22335
rect 29771 22272 29837 22275
rect 30105 22270 30175 22275
rect 30376 22306 30446 22311
rect 31887 22306 31953 22309
rect 30376 22246 30381 22306
rect 30441 22304 31953 22306
rect 30441 22248 31892 22304
rect 31948 22248 31953 22304
rect 30441 22246 31953 22248
rect 30376 22241 30446 22246
rect 31887 22243 31953 22246
rect 15256 4203 15322 4206
rect 19925 4203 19995 4208
rect 15256 4201 19930 4203
rect 15256 4145 15261 4201
rect 15317 4145 19930 4201
rect 15256 4143 19930 4145
rect 19990 4143 19995 4203
rect 15256 4140 15322 4143
rect 19925 4138 19995 4143
rect 18491 3531 18561 3536
rect 19681 3531 19747 3534
rect 18491 3471 18496 3531
rect 18556 3529 19747 3531
rect 18556 3473 19686 3529
rect 19742 3473 19747 3529
rect 18556 3471 19747 3473
rect 18491 3466 18561 3471
rect 19681 3468 19747 3471
<< via3 >>
rect -38 75288 350 75676
rect 44459 75288 44847 75676
rect 422 74828 810 75216
rect 43999 74828 44387 75216
rect 882 74368 1270 74756
rect 43539 74368 43927 74756
rect 1342 73908 1730 74296
rect 43079 73908 43467 74296
rect 1342 45799 1730 46187
rect 43079 45799 43467 46187
rect 882 45339 1270 45727
rect 43539 45339 43927 45727
rect 422 44879 810 45267
rect 43999 44879 44387 45267
rect -38 44419 350 44807
rect 44459 44419 44847 44807
<< metal4 >>
rect -44 75676 356 75683
rect -44 75288 -38 75676
rect 350 75288 356 75676
rect -44 44807 356 75288
rect -44 44419 -38 44807
rect 350 44419 356 44807
rect -44 44413 356 44419
rect 416 75216 816 75683
rect 416 74828 422 75216
rect 810 74828 816 75216
rect 416 45267 816 74828
rect 416 44879 422 45267
rect 810 44879 816 45267
rect 416 44413 816 44879
rect 876 74756 1276 75683
rect 876 74368 882 74756
rect 1270 74368 1276 74756
rect 876 45727 1276 74368
rect 876 45339 882 45727
rect 1270 45339 1276 45727
rect 876 44413 1276 45339
rect 1336 74296 1736 75683
rect 1336 73908 1342 74296
rect 1730 73908 1736 74296
rect 1336 54039 1736 73908
rect 43073 74296 43473 75683
rect 43073 73908 43079 74296
rect 43467 73908 43473 74296
rect 1336 53637 1740 54039
rect 1336 46187 1736 53637
rect 1336 45799 1342 46187
rect 1730 45799 1736 46187
rect 1336 44413 1736 45799
rect 43073 46187 43473 73908
rect 43073 45799 43079 46187
rect 43467 45799 43473 46187
rect 43073 44413 43473 45799
rect 43533 74756 43933 75683
rect 43533 74368 43539 74756
rect 43927 74368 43933 74756
rect 43533 45727 43933 74368
rect 43533 45339 43539 45727
rect 43927 45339 43933 45727
rect 43533 44413 43933 45339
rect 43993 75216 44393 75683
rect 43993 74828 43999 75216
rect 44387 74828 44393 75216
rect 43993 45267 44393 74828
rect 43993 44879 43999 45267
rect 44387 44879 44393 45267
rect 43993 44413 44393 44879
rect 44453 75676 44853 75683
rect 44453 75288 44459 75676
rect 44847 75288 44853 75676
rect 44453 44807 44853 75288
rect 44453 44419 44459 44807
rect 44847 44419 44853 44807
rect 44453 44413 44853 44419
use brownout_ana  brownout_ana_0 ~/chipalooza/sky130_ajc_ip__brownout/mag
timestamp 1712901199
transform 1 0 29373 0 1 25849
box -29373 -25849 12300 13900
use brownout_dig  brownout_dig_0
timestamp 1712897939
transform 1 0 30384 0 1 26140
box 0 0 11173 13317
<< labels >>
flabel metal3 3283 44873 3283 44873 0 FreeSans 1600 0 0 0 dvss
port 4 nsew
flabel metal3 3283 45333 3283 45333 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 3283 45793 3283 45793 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal3 3283 44413 3283 44413 0 FreeSans 1600 0 0 0 dvdd
port 3 nsew
<< end >>

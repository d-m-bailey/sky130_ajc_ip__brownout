magic
tech sky130A
magscale 1 2
timestamp 1712930986
<< nwell >>
rect -5203 -1457 5203 1457
<< mvpmos >>
rect -4945 1030 -3345 1230
rect -3287 1030 -1687 1230
rect -1629 1030 -29 1230
rect 29 1030 1629 1230
rect 1687 1030 3287 1230
rect 3345 1030 4945 1230
rect -4945 665 -3345 865
rect -3287 665 -1687 865
rect -1629 665 -29 865
rect 29 665 1629 865
rect 1687 665 3287 865
rect 3345 665 4945 865
rect -4945 300 -3345 500
rect -3287 300 -1687 500
rect -1629 300 -29 500
rect 29 300 1629 500
rect 1687 300 3287 500
rect 3345 300 4945 500
rect -4945 -65 -3345 135
rect -3287 -65 -1687 135
rect -1629 -65 -29 135
rect 29 -65 1629 135
rect 1687 -65 3287 135
rect 3345 -65 4945 135
rect -4945 -430 -3345 -230
rect -3287 -430 -1687 -230
rect -1629 -430 -29 -230
rect 29 -430 1629 -230
rect 1687 -430 3287 -230
rect 3345 -430 4945 -230
rect -4945 -795 -3345 -595
rect -3287 -795 -1687 -595
rect -1629 -795 -29 -595
rect 29 -795 1629 -595
rect 1687 -795 3287 -595
rect 3345 -795 4945 -595
rect -4945 -1160 -3345 -960
rect -3287 -1160 -1687 -960
rect -1629 -1160 -29 -960
rect 29 -1160 1629 -960
rect 1687 -1160 3287 -960
rect 3345 -1160 4945 -960
<< mvpdiff >>
rect -5003 1218 -4945 1230
rect -5003 1042 -4991 1218
rect -4957 1042 -4945 1218
rect -5003 1030 -4945 1042
rect -3345 1218 -3287 1230
rect -3345 1042 -3333 1218
rect -3299 1042 -3287 1218
rect -3345 1030 -3287 1042
rect -1687 1218 -1629 1230
rect -1687 1042 -1675 1218
rect -1641 1042 -1629 1218
rect -1687 1030 -1629 1042
rect -29 1218 29 1230
rect -29 1042 -17 1218
rect 17 1042 29 1218
rect -29 1030 29 1042
rect 1629 1218 1687 1230
rect 1629 1042 1641 1218
rect 1675 1042 1687 1218
rect 1629 1030 1687 1042
rect 3287 1218 3345 1230
rect 3287 1042 3299 1218
rect 3333 1042 3345 1218
rect 3287 1030 3345 1042
rect 4945 1218 5003 1230
rect 4945 1042 4957 1218
rect 4991 1042 5003 1218
rect 4945 1030 5003 1042
rect -5003 853 -4945 865
rect -5003 677 -4991 853
rect -4957 677 -4945 853
rect -5003 665 -4945 677
rect -3345 853 -3287 865
rect -3345 677 -3333 853
rect -3299 677 -3287 853
rect -3345 665 -3287 677
rect -1687 853 -1629 865
rect -1687 677 -1675 853
rect -1641 677 -1629 853
rect -1687 665 -1629 677
rect -29 853 29 865
rect -29 677 -17 853
rect 17 677 29 853
rect -29 665 29 677
rect 1629 853 1687 865
rect 1629 677 1641 853
rect 1675 677 1687 853
rect 1629 665 1687 677
rect 3287 853 3345 865
rect 3287 677 3299 853
rect 3333 677 3345 853
rect 3287 665 3345 677
rect 4945 853 5003 865
rect 4945 677 4957 853
rect 4991 677 5003 853
rect 4945 665 5003 677
rect -5003 488 -4945 500
rect -5003 312 -4991 488
rect -4957 312 -4945 488
rect -5003 300 -4945 312
rect -3345 488 -3287 500
rect -3345 312 -3333 488
rect -3299 312 -3287 488
rect -3345 300 -3287 312
rect -1687 488 -1629 500
rect -1687 312 -1675 488
rect -1641 312 -1629 488
rect -1687 300 -1629 312
rect -29 488 29 500
rect -29 312 -17 488
rect 17 312 29 488
rect -29 300 29 312
rect 1629 488 1687 500
rect 1629 312 1641 488
rect 1675 312 1687 488
rect 1629 300 1687 312
rect 3287 488 3345 500
rect 3287 312 3299 488
rect 3333 312 3345 488
rect 3287 300 3345 312
rect 4945 488 5003 500
rect 4945 312 4957 488
rect 4991 312 5003 488
rect 4945 300 5003 312
rect -5003 123 -4945 135
rect -5003 -53 -4991 123
rect -4957 -53 -4945 123
rect -5003 -65 -4945 -53
rect -3345 123 -3287 135
rect -3345 -53 -3333 123
rect -3299 -53 -3287 123
rect -3345 -65 -3287 -53
rect -1687 123 -1629 135
rect -1687 -53 -1675 123
rect -1641 -53 -1629 123
rect -1687 -65 -1629 -53
rect -29 123 29 135
rect -29 -53 -17 123
rect 17 -53 29 123
rect -29 -65 29 -53
rect 1629 123 1687 135
rect 1629 -53 1641 123
rect 1675 -53 1687 123
rect 1629 -65 1687 -53
rect 3287 123 3345 135
rect 3287 -53 3299 123
rect 3333 -53 3345 123
rect 3287 -65 3345 -53
rect 4945 123 5003 135
rect 4945 -53 4957 123
rect 4991 -53 5003 123
rect 4945 -65 5003 -53
rect -5003 -242 -4945 -230
rect -5003 -418 -4991 -242
rect -4957 -418 -4945 -242
rect -5003 -430 -4945 -418
rect -3345 -242 -3287 -230
rect -3345 -418 -3333 -242
rect -3299 -418 -3287 -242
rect -3345 -430 -3287 -418
rect -1687 -242 -1629 -230
rect -1687 -418 -1675 -242
rect -1641 -418 -1629 -242
rect -1687 -430 -1629 -418
rect -29 -242 29 -230
rect -29 -418 -17 -242
rect 17 -418 29 -242
rect -29 -430 29 -418
rect 1629 -242 1687 -230
rect 1629 -418 1641 -242
rect 1675 -418 1687 -242
rect 1629 -430 1687 -418
rect 3287 -242 3345 -230
rect 3287 -418 3299 -242
rect 3333 -418 3345 -242
rect 3287 -430 3345 -418
rect 4945 -242 5003 -230
rect 4945 -418 4957 -242
rect 4991 -418 5003 -242
rect 4945 -430 5003 -418
rect -5003 -607 -4945 -595
rect -5003 -783 -4991 -607
rect -4957 -783 -4945 -607
rect -5003 -795 -4945 -783
rect -3345 -607 -3287 -595
rect -3345 -783 -3333 -607
rect -3299 -783 -3287 -607
rect -3345 -795 -3287 -783
rect -1687 -607 -1629 -595
rect -1687 -783 -1675 -607
rect -1641 -783 -1629 -607
rect -1687 -795 -1629 -783
rect -29 -607 29 -595
rect -29 -783 -17 -607
rect 17 -783 29 -607
rect -29 -795 29 -783
rect 1629 -607 1687 -595
rect 1629 -783 1641 -607
rect 1675 -783 1687 -607
rect 1629 -795 1687 -783
rect 3287 -607 3345 -595
rect 3287 -783 3299 -607
rect 3333 -783 3345 -607
rect 3287 -795 3345 -783
rect 4945 -607 5003 -595
rect 4945 -783 4957 -607
rect 4991 -783 5003 -607
rect 4945 -795 5003 -783
rect -5003 -972 -4945 -960
rect -5003 -1148 -4991 -972
rect -4957 -1148 -4945 -972
rect -5003 -1160 -4945 -1148
rect -3345 -972 -3287 -960
rect -3345 -1148 -3333 -972
rect -3299 -1148 -3287 -972
rect -3345 -1160 -3287 -1148
rect -1687 -972 -1629 -960
rect -1687 -1148 -1675 -972
rect -1641 -1148 -1629 -972
rect -1687 -1160 -1629 -1148
rect -29 -972 29 -960
rect -29 -1148 -17 -972
rect 17 -1148 29 -972
rect -29 -1160 29 -1148
rect 1629 -972 1687 -960
rect 1629 -1148 1641 -972
rect 1675 -1148 1687 -972
rect 1629 -1160 1687 -1148
rect 3287 -972 3345 -960
rect 3287 -1148 3299 -972
rect 3333 -1148 3345 -972
rect 3287 -1160 3345 -1148
rect 4945 -972 5003 -960
rect 4945 -1148 4957 -972
rect 4991 -1148 5003 -972
rect 4945 -1160 5003 -1148
<< mvpdiffc >>
rect -4991 1042 -4957 1218
rect -3333 1042 -3299 1218
rect -1675 1042 -1641 1218
rect -17 1042 17 1218
rect 1641 1042 1675 1218
rect 3299 1042 3333 1218
rect 4957 1042 4991 1218
rect -4991 677 -4957 853
rect -3333 677 -3299 853
rect -1675 677 -1641 853
rect -17 677 17 853
rect 1641 677 1675 853
rect 3299 677 3333 853
rect 4957 677 4991 853
rect -4991 312 -4957 488
rect -3333 312 -3299 488
rect -1675 312 -1641 488
rect -17 312 17 488
rect 1641 312 1675 488
rect 3299 312 3333 488
rect 4957 312 4991 488
rect -4991 -53 -4957 123
rect -3333 -53 -3299 123
rect -1675 -53 -1641 123
rect -17 -53 17 123
rect 1641 -53 1675 123
rect 3299 -53 3333 123
rect 4957 -53 4991 123
rect -4991 -418 -4957 -242
rect -3333 -418 -3299 -242
rect -1675 -418 -1641 -242
rect -17 -418 17 -242
rect 1641 -418 1675 -242
rect 3299 -418 3333 -242
rect 4957 -418 4991 -242
rect -4991 -783 -4957 -607
rect -3333 -783 -3299 -607
rect -1675 -783 -1641 -607
rect -17 -783 17 -607
rect 1641 -783 1675 -607
rect 3299 -783 3333 -607
rect 4957 -783 4991 -607
rect -4991 -1148 -4957 -972
rect -3333 -1148 -3299 -972
rect -1675 -1148 -1641 -972
rect -17 -1148 17 -972
rect 1641 -1148 1675 -972
rect 3299 -1148 3333 -972
rect 4957 -1148 4991 -972
<< mvnsubdiff >>
rect -5137 1379 5137 1391
rect -5137 1345 -5029 1379
rect 5029 1345 5137 1379
rect -5137 1333 5137 1345
rect -5137 1283 -5079 1333
rect -5137 -1283 -5125 1283
rect -5091 -1283 -5079 1283
rect 5079 1283 5137 1333
rect -5137 -1333 -5079 -1283
rect 5079 -1283 5091 1283
rect 5125 -1283 5137 1283
rect 5079 -1333 5137 -1283
rect -5137 -1345 5137 -1333
rect -5137 -1379 -5029 -1345
rect 5029 -1379 5137 -1345
rect -5137 -1391 5137 -1379
<< mvnsubdiffcont >>
rect -5029 1345 5029 1379
rect -5125 -1283 -5091 1283
rect 5091 -1283 5125 1283
rect -5029 -1379 5029 -1345
<< poly >>
rect -4945 1230 -3345 1256
rect -3287 1230 -1687 1256
rect -1629 1230 -29 1256
rect 29 1230 1629 1256
rect 1687 1230 3287 1256
rect 3345 1230 4945 1256
rect -4945 983 -3345 1030
rect -4945 949 -4929 983
rect -3361 949 -3345 983
rect -4945 933 -3345 949
rect -3287 983 -1687 1030
rect -3287 949 -3271 983
rect -1703 949 -1687 983
rect -3287 933 -1687 949
rect -1629 983 -29 1030
rect -1629 949 -1613 983
rect -45 949 -29 983
rect -1629 933 -29 949
rect 29 983 1629 1030
rect 29 949 45 983
rect 1613 949 1629 983
rect 29 933 1629 949
rect 1687 983 3287 1030
rect 1687 949 1703 983
rect 3271 949 3287 983
rect 1687 933 3287 949
rect 3345 983 4945 1030
rect 3345 949 3361 983
rect 4929 949 4945 983
rect 3345 933 4945 949
rect -4945 865 -3345 891
rect -3287 865 -1687 891
rect -1629 865 -29 891
rect 29 865 1629 891
rect 1687 865 3287 891
rect 3345 865 4945 891
rect -4945 618 -3345 665
rect -4945 584 -4929 618
rect -3361 584 -3345 618
rect -4945 568 -3345 584
rect -3287 618 -1687 665
rect -3287 584 -3271 618
rect -1703 584 -1687 618
rect -3287 568 -1687 584
rect -1629 618 -29 665
rect -1629 584 -1613 618
rect -45 584 -29 618
rect -1629 568 -29 584
rect 29 618 1629 665
rect 29 584 45 618
rect 1613 584 1629 618
rect 29 568 1629 584
rect 1687 618 3287 665
rect 1687 584 1703 618
rect 3271 584 3287 618
rect 1687 568 3287 584
rect 3345 618 4945 665
rect 3345 584 3361 618
rect 4929 584 4945 618
rect 3345 568 4945 584
rect -4945 500 -3345 526
rect -3287 500 -1687 526
rect -1629 500 -29 526
rect 29 500 1629 526
rect 1687 500 3287 526
rect 3345 500 4945 526
rect -4945 253 -3345 300
rect -4945 219 -4929 253
rect -3361 219 -3345 253
rect -4945 203 -3345 219
rect -3287 253 -1687 300
rect -3287 219 -3271 253
rect -1703 219 -1687 253
rect -3287 203 -1687 219
rect -1629 253 -29 300
rect -1629 219 -1613 253
rect -45 219 -29 253
rect -1629 203 -29 219
rect 29 253 1629 300
rect 29 219 45 253
rect 1613 219 1629 253
rect 29 203 1629 219
rect 1687 253 3287 300
rect 1687 219 1703 253
rect 3271 219 3287 253
rect 1687 203 3287 219
rect 3345 253 4945 300
rect 3345 219 3361 253
rect 4929 219 4945 253
rect 3345 203 4945 219
rect -4945 135 -3345 161
rect -3287 135 -1687 161
rect -1629 135 -29 161
rect 29 135 1629 161
rect 1687 135 3287 161
rect 3345 135 4945 161
rect -4945 -112 -3345 -65
rect -4945 -146 -4929 -112
rect -3361 -146 -3345 -112
rect -4945 -162 -3345 -146
rect -3287 -112 -1687 -65
rect -3287 -146 -3271 -112
rect -1703 -146 -1687 -112
rect -3287 -162 -1687 -146
rect -1629 -112 -29 -65
rect -1629 -146 -1613 -112
rect -45 -146 -29 -112
rect -1629 -162 -29 -146
rect 29 -112 1629 -65
rect 29 -146 45 -112
rect 1613 -146 1629 -112
rect 29 -162 1629 -146
rect 1687 -112 3287 -65
rect 1687 -146 1703 -112
rect 3271 -146 3287 -112
rect 1687 -162 3287 -146
rect 3345 -112 4945 -65
rect 3345 -146 3361 -112
rect 4929 -146 4945 -112
rect 3345 -162 4945 -146
rect -4945 -230 -3345 -204
rect -3287 -230 -1687 -204
rect -1629 -230 -29 -204
rect 29 -230 1629 -204
rect 1687 -230 3287 -204
rect 3345 -230 4945 -204
rect -4945 -477 -3345 -430
rect -4945 -511 -4929 -477
rect -3361 -511 -3345 -477
rect -4945 -527 -3345 -511
rect -3287 -477 -1687 -430
rect -3287 -511 -3271 -477
rect -1703 -511 -1687 -477
rect -3287 -527 -1687 -511
rect -1629 -477 -29 -430
rect -1629 -511 -1613 -477
rect -45 -511 -29 -477
rect -1629 -527 -29 -511
rect 29 -477 1629 -430
rect 29 -511 45 -477
rect 1613 -511 1629 -477
rect 29 -527 1629 -511
rect 1687 -477 3287 -430
rect 1687 -511 1703 -477
rect 3271 -511 3287 -477
rect 1687 -527 3287 -511
rect 3345 -477 4945 -430
rect 3345 -511 3361 -477
rect 4929 -511 4945 -477
rect 3345 -527 4945 -511
rect -4945 -595 -3345 -569
rect -3287 -595 -1687 -569
rect -1629 -595 -29 -569
rect 29 -595 1629 -569
rect 1687 -595 3287 -569
rect 3345 -595 4945 -569
rect -4945 -842 -3345 -795
rect -4945 -876 -4929 -842
rect -3361 -876 -3345 -842
rect -4945 -892 -3345 -876
rect -3287 -842 -1687 -795
rect -3287 -876 -3271 -842
rect -1703 -876 -1687 -842
rect -3287 -892 -1687 -876
rect -1629 -842 -29 -795
rect -1629 -876 -1613 -842
rect -45 -876 -29 -842
rect -1629 -892 -29 -876
rect 29 -842 1629 -795
rect 29 -876 45 -842
rect 1613 -876 1629 -842
rect 29 -892 1629 -876
rect 1687 -842 3287 -795
rect 1687 -876 1703 -842
rect 3271 -876 3287 -842
rect 1687 -892 3287 -876
rect 3345 -842 4945 -795
rect 3345 -876 3361 -842
rect 4929 -876 4945 -842
rect 3345 -892 4945 -876
rect -4945 -960 -3345 -934
rect -3287 -960 -1687 -934
rect -1629 -960 -29 -934
rect 29 -960 1629 -934
rect 1687 -960 3287 -934
rect 3345 -960 4945 -934
rect -4945 -1207 -3345 -1160
rect -4945 -1241 -4929 -1207
rect -3361 -1241 -3345 -1207
rect -4945 -1257 -3345 -1241
rect -3287 -1207 -1687 -1160
rect -3287 -1241 -3271 -1207
rect -1703 -1241 -1687 -1207
rect -3287 -1257 -1687 -1241
rect -1629 -1207 -29 -1160
rect -1629 -1241 -1613 -1207
rect -45 -1241 -29 -1207
rect -1629 -1257 -29 -1241
rect 29 -1207 1629 -1160
rect 29 -1241 45 -1207
rect 1613 -1241 1629 -1207
rect 29 -1257 1629 -1241
rect 1687 -1207 3287 -1160
rect 1687 -1241 1703 -1207
rect 3271 -1241 3287 -1207
rect 1687 -1257 3287 -1241
rect 3345 -1207 4945 -1160
rect 3345 -1241 3361 -1207
rect 4929 -1241 4945 -1207
rect 3345 -1257 4945 -1241
<< polycont >>
rect -4929 949 -3361 983
rect -3271 949 -1703 983
rect -1613 949 -45 983
rect 45 949 1613 983
rect 1703 949 3271 983
rect 3361 949 4929 983
rect -4929 584 -3361 618
rect -3271 584 -1703 618
rect -1613 584 -45 618
rect 45 584 1613 618
rect 1703 584 3271 618
rect 3361 584 4929 618
rect -4929 219 -3361 253
rect -3271 219 -1703 253
rect -1613 219 -45 253
rect 45 219 1613 253
rect 1703 219 3271 253
rect 3361 219 4929 253
rect -4929 -146 -3361 -112
rect -3271 -146 -1703 -112
rect -1613 -146 -45 -112
rect 45 -146 1613 -112
rect 1703 -146 3271 -112
rect 3361 -146 4929 -112
rect -4929 -511 -3361 -477
rect -3271 -511 -1703 -477
rect -1613 -511 -45 -477
rect 45 -511 1613 -477
rect 1703 -511 3271 -477
rect 3361 -511 4929 -477
rect -4929 -876 -3361 -842
rect -3271 -876 -1703 -842
rect -1613 -876 -45 -842
rect 45 -876 1613 -842
rect 1703 -876 3271 -842
rect 3361 -876 4929 -842
rect -4929 -1241 -3361 -1207
rect -3271 -1241 -1703 -1207
rect -1613 -1241 -45 -1207
rect 45 -1241 1613 -1207
rect 1703 -1241 3271 -1207
rect 3361 -1241 4929 -1207
<< locali >>
rect -5125 1345 -5029 1379
rect 5029 1345 5125 1379
rect -5125 1283 -5091 1345
rect 5091 1283 5125 1345
rect -4991 1218 -4957 1234
rect -4991 1026 -4957 1042
rect -3333 1218 -3299 1234
rect -3333 1026 -3299 1042
rect -1675 1218 -1641 1234
rect -1675 1026 -1641 1042
rect -17 1218 17 1234
rect -17 1026 17 1042
rect 1641 1218 1675 1234
rect 1641 1026 1675 1042
rect 3299 1218 3333 1234
rect 3299 1026 3333 1042
rect 4957 1218 4991 1234
rect 4957 1026 4991 1042
rect -4945 949 -4929 983
rect -3361 949 -3345 983
rect -3287 949 -3271 983
rect -1703 949 -1687 983
rect -1629 949 -1613 983
rect -45 949 -29 983
rect 29 949 45 983
rect 1613 949 1629 983
rect 1687 949 1703 983
rect 3271 949 3287 983
rect 3345 949 3361 983
rect 4929 949 4945 983
rect -4991 853 -4957 869
rect -4991 661 -4957 677
rect -3333 853 -3299 869
rect -3333 661 -3299 677
rect -1675 853 -1641 869
rect -1675 661 -1641 677
rect -17 853 17 869
rect -17 661 17 677
rect 1641 853 1675 869
rect 1641 661 1675 677
rect 3299 853 3333 869
rect 3299 661 3333 677
rect 4957 853 4991 869
rect 4957 661 4991 677
rect -4945 584 -4929 618
rect -3361 584 -3345 618
rect -3287 584 -3271 618
rect -1703 584 -1687 618
rect -1629 584 -1613 618
rect -45 584 -29 618
rect 29 584 45 618
rect 1613 584 1629 618
rect 1687 584 1703 618
rect 3271 584 3287 618
rect 3345 584 3361 618
rect 4929 584 4945 618
rect -4991 488 -4957 504
rect -4991 296 -4957 312
rect -3333 488 -3299 504
rect -3333 296 -3299 312
rect -1675 488 -1641 504
rect -1675 296 -1641 312
rect -17 488 17 504
rect -17 296 17 312
rect 1641 488 1675 504
rect 1641 296 1675 312
rect 3299 488 3333 504
rect 3299 296 3333 312
rect 4957 488 4991 504
rect 4957 296 4991 312
rect -4945 219 -4929 253
rect -3361 219 -3345 253
rect -3287 219 -3271 253
rect -1703 219 -1687 253
rect -1629 219 -1613 253
rect -45 219 -29 253
rect 29 219 45 253
rect 1613 219 1629 253
rect 1687 219 1703 253
rect 3271 219 3287 253
rect 3345 219 3361 253
rect 4929 219 4945 253
rect -4991 123 -4957 139
rect -4991 -69 -4957 -53
rect -3333 123 -3299 139
rect -3333 -69 -3299 -53
rect -1675 123 -1641 139
rect -1675 -69 -1641 -53
rect -17 123 17 139
rect -17 -69 17 -53
rect 1641 123 1675 139
rect 1641 -69 1675 -53
rect 3299 123 3333 139
rect 3299 -69 3333 -53
rect 4957 123 4991 139
rect 4957 -69 4991 -53
rect -4945 -146 -4929 -112
rect -3361 -146 -3345 -112
rect -3287 -146 -3271 -112
rect -1703 -146 -1687 -112
rect -1629 -146 -1613 -112
rect -45 -146 -29 -112
rect 29 -146 45 -112
rect 1613 -146 1629 -112
rect 1687 -146 1703 -112
rect 3271 -146 3287 -112
rect 3345 -146 3361 -112
rect 4929 -146 4945 -112
rect -4991 -242 -4957 -226
rect -4991 -434 -4957 -418
rect -3333 -242 -3299 -226
rect -3333 -434 -3299 -418
rect -1675 -242 -1641 -226
rect -1675 -434 -1641 -418
rect -17 -242 17 -226
rect -17 -434 17 -418
rect 1641 -242 1675 -226
rect 1641 -434 1675 -418
rect 3299 -242 3333 -226
rect 3299 -434 3333 -418
rect 4957 -242 4991 -226
rect 4957 -434 4991 -418
rect -4945 -511 -4929 -477
rect -3361 -511 -3345 -477
rect -3287 -511 -3271 -477
rect -1703 -511 -1687 -477
rect -1629 -511 -1613 -477
rect -45 -511 -29 -477
rect 29 -511 45 -477
rect 1613 -511 1629 -477
rect 1687 -511 1703 -477
rect 3271 -511 3287 -477
rect 3345 -511 3361 -477
rect 4929 -511 4945 -477
rect -4991 -607 -4957 -591
rect -4991 -799 -4957 -783
rect -3333 -607 -3299 -591
rect -3333 -799 -3299 -783
rect -1675 -607 -1641 -591
rect -1675 -799 -1641 -783
rect -17 -607 17 -591
rect -17 -799 17 -783
rect 1641 -607 1675 -591
rect 1641 -799 1675 -783
rect 3299 -607 3333 -591
rect 3299 -799 3333 -783
rect 4957 -607 4991 -591
rect 4957 -799 4991 -783
rect -4945 -876 -4929 -842
rect -3361 -876 -3345 -842
rect -3287 -876 -3271 -842
rect -1703 -876 -1687 -842
rect -1629 -876 -1613 -842
rect -45 -876 -29 -842
rect 29 -876 45 -842
rect 1613 -876 1629 -842
rect 1687 -876 1703 -842
rect 3271 -876 3287 -842
rect 3345 -876 3361 -842
rect 4929 -876 4945 -842
rect -4991 -972 -4957 -956
rect -4991 -1164 -4957 -1148
rect -3333 -972 -3299 -956
rect -3333 -1164 -3299 -1148
rect -1675 -972 -1641 -956
rect -1675 -1164 -1641 -1148
rect -17 -972 17 -956
rect -17 -1164 17 -1148
rect 1641 -972 1675 -956
rect 1641 -1164 1675 -1148
rect 3299 -972 3333 -956
rect 3299 -1164 3333 -1148
rect 4957 -972 4991 -956
rect 4957 -1164 4991 -1148
rect -4945 -1241 -4929 -1207
rect -3361 -1241 -3345 -1207
rect -3287 -1241 -3271 -1207
rect -1703 -1241 -1687 -1207
rect -1629 -1241 -1613 -1207
rect -45 -1241 -29 -1207
rect 29 -1241 45 -1207
rect 1613 -1241 1629 -1207
rect 1687 -1241 1703 -1207
rect 3271 -1241 3287 -1207
rect 3345 -1241 3361 -1207
rect 4929 -1241 4945 -1207
rect -5125 -1345 -5091 -1283
rect 5091 -1345 5125 -1283
rect -5125 -1379 -5029 -1345
rect 5029 -1379 5125 -1345
<< viali >>
rect -4991 1042 -4957 1218
rect -3333 1042 -3299 1218
rect -1675 1042 -1641 1218
rect -17 1042 17 1218
rect 1641 1042 1675 1218
rect 3299 1042 3333 1218
rect 4957 1042 4991 1218
rect -4929 949 -3361 983
rect -3271 949 -1703 983
rect -1613 949 -45 983
rect 45 949 1613 983
rect 1703 949 3271 983
rect 3361 949 4929 983
rect -4991 677 -4957 853
rect -3333 677 -3299 853
rect -1675 677 -1641 853
rect -17 677 17 853
rect 1641 677 1675 853
rect 3299 677 3333 853
rect 4957 677 4991 853
rect -4929 584 -3361 618
rect -3271 584 -1703 618
rect -1613 584 -45 618
rect 45 584 1613 618
rect 1703 584 3271 618
rect 3361 584 4929 618
rect -4991 312 -4957 488
rect -3333 312 -3299 488
rect -1675 312 -1641 488
rect -17 312 17 488
rect 1641 312 1675 488
rect 3299 312 3333 488
rect 4957 312 4991 488
rect -4929 219 -3361 253
rect -3271 219 -1703 253
rect -1613 219 -45 253
rect 45 219 1613 253
rect 1703 219 3271 253
rect 3361 219 4929 253
rect -4991 -53 -4957 123
rect -3333 -53 -3299 123
rect -1675 -53 -1641 123
rect -17 -53 17 123
rect 1641 -53 1675 123
rect 3299 -53 3333 123
rect 4957 -53 4991 123
rect -4929 -146 -3361 -112
rect -3271 -146 -1703 -112
rect -1613 -146 -45 -112
rect 45 -146 1613 -112
rect 1703 -146 3271 -112
rect 3361 -146 4929 -112
rect -4991 -418 -4957 -242
rect -3333 -418 -3299 -242
rect -1675 -418 -1641 -242
rect -17 -418 17 -242
rect 1641 -418 1675 -242
rect 3299 -418 3333 -242
rect 4957 -418 4991 -242
rect -4929 -511 -3361 -477
rect -3271 -511 -1703 -477
rect -1613 -511 -45 -477
rect 45 -511 1613 -477
rect 1703 -511 3271 -477
rect 3361 -511 4929 -477
rect -4991 -783 -4957 -607
rect -3333 -783 -3299 -607
rect -1675 -783 -1641 -607
rect -17 -783 17 -607
rect 1641 -783 1675 -607
rect 3299 -783 3333 -607
rect 4957 -783 4991 -607
rect -4929 -876 -3361 -842
rect -3271 -876 -1703 -842
rect -1613 -876 -45 -842
rect 45 -876 1613 -842
rect 1703 -876 3271 -842
rect 3361 -876 4929 -842
rect -4991 -1148 -4957 -972
rect -3333 -1148 -3299 -972
rect -1675 -1148 -1641 -972
rect -17 -1148 17 -972
rect 1641 -1148 1675 -972
rect 3299 -1148 3333 -972
rect 4957 -1148 4991 -972
rect -4929 -1241 -3361 -1207
rect -3271 -1241 -1703 -1207
rect -1613 -1241 -45 -1207
rect 45 -1241 1613 -1207
rect 1703 -1241 3271 -1207
rect 3361 -1241 4929 -1207
<< metal1 >>
rect -4997 1218 -4951 1230
rect -4997 1042 -4991 1218
rect -4957 1042 -4951 1218
rect -4997 1030 -4951 1042
rect -3339 1218 -3293 1230
rect -3339 1042 -3333 1218
rect -3299 1042 -3293 1218
rect -3339 1030 -3293 1042
rect -1681 1218 -1635 1230
rect -1681 1042 -1675 1218
rect -1641 1042 -1635 1218
rect -1681 1030 -1635 1042
rect -23 1218 23 1230
rect -23 1042 -17 1218
rect 17 1042 23 1218
rect -23 1030 23 1042
rect 1635 1218 1681 1230
rect 1635 1042 1641 1218
rect 1675 1042 1681 1218
rect 1635 1030 1681 1042
rect 3293 1218 3339 1230
rect 3293 1042 3299 1218
rect 3333 1042 3339 1218
rect 3293 1030 3339 1042
rect 4951 1218 4997 1230
rect 4951 1042 4957 1218
rect 4991 1042 4997 1218
rect 4951 1030 4997 1042
rect -4941 983 -3349 989
rect -4941 949 -4929 983
rect -3361 949 -3349 983
rect -4941 943 -3349 949
rect -3283 983 -1691 989
rect -3283 949 -3271 983
rect -1703 949 -1691 983
rect -3283 943 -1691 949
rect -1625 983 -33 989
rect -1625 949 -1613 983
rect -45 949 -33 983
rect -1625 943 -33 949
rect 33 983 1625 989
rect 33 949 45 983
rect 1613 949 1625 983
rect 33 943 1625 949
rect 1691 983 3283 989
rect 1691 949 1703 983
rect 3271 949 3283 983
rect 1691 943 3283 949
rect 3349 983 4941 989
rect 3349 949 3361 983
rect 4929 949 4941 983
rect 3349 943 4941 949
rect -4997 853 -4951 865
rect -4997 677 -4991 853
rect -4957 677 -4951 853
rect -4997 665 -4951 677
rect -3339 853 -3293 865
rect -3339 677 -3333 853
rect -3299 677 -3293 853
rect -3339 665 -3293 677
rect -1681 853 -1635 865
rect -1681 677 -1675 853
rect -1641 677 -1635 853
rect -1681 665 -1635 677
rect -23 853 23 865
rect -23 677 -17 853
rect 17 677 23 853
rect -23 665 23 677
rect 1635 853 1681 865
rect 1635 677 1641 853
rect 1675 677 1681 853
rect 1635 665 1681 677
rect 3293 853 3339 865
rect 3293 677 3299 853
rect 3333 677 3339 853
rect 3293 665 3339 677
rect 4951 853 4997 865
rect 4951 677 4957 853
rect 4991 677 4997 853
rect 4951 665 4997 677
rect -4941 618 -3349 624
rect -4941 584 -4929 618
rect -3361 584 -3349 618
rect -4941 578 -3349 584
rect -3283 618 -1691 624
rect -3283 584 -3271 618
rect -1703 584 -1691 618
rect -3283 578 -1691 584
rect -1625 618 -33 624
rect -1625 584 -1613 618
rect -45 584 -33 618
rect -1625 578 -33 584
rect 33 618 1625 624
rect 33 584 45 618
rect 1613 584 1625 618
rect 33 578 1625 584
rect 1691 618 3283 624
rect 1691 584 1703 618
rect 3271 584 3283 618
rect 1691 578 3283 584
rect 3349 618 4941 624
rect 3349 584 3361 618
rect 4929 584 4941 618
rect 3349 578 4941 584
rect -4997 488 -4951 500
rect -4997 312 -4991 488
rect -4957 312 -4951 488
rect -4997 300 -4951 312
rect -3339 488 -3293 500
rect -3339 312 -3333 488
rect -3299 312 -3293 488
rect -3339 300 -3293 312
rect -1681 488 -1635 500
rect -1681 312 -1675 488
rect -1641 312 -1635 488
rect -1681 300 -1635 312
rect -23 488 23 500
rect -23 312 -17 488
rect 17 312 23 488
rect -23 300 23 312
rect 1635 488 1681 500
rect 1635 312 1641 488
rect 1675 312 1681 488
rect 1635 300 1681 312
rect 3293 488 3339 500
rect 3293 312 3299 488
rect 3333 312 3339 488
rect 3293 300 3339 312
rect 4951 488 4997 500
rect 4951 312 4957 488
rect 4991 312 4997 488
rect 4951 300 4997 312
rect -4941 253 -3349 259
rect -4941 219 -4929 253
rect -3361 219 -3349 253
rect -4941 213 -3349 219
rect -3283 253 -1691 259
rect -3283 219 -3271 253
rect -1703 219 -1691 253
rect -3283 213 -1691 219
rect -1625 253 -33 259
rect -1625 219 -1613 253
rect -45 219 -33 253
rect -1625 213 -33 219
rect 33 253 1625 259
rect 33 219 45 253
rect 1613 219 1625 253
rect 33 213 1625 219
rect 1691 253 3283 259
rect 1691 219 1703 253
rect 3271 219 3283 253
rect 1691 213 3283 219
rect 3349 253 4941 259
rect 3349 219 3361 253
rect 4929 219 4941 253
rect 3349 213 4941 219
rect -4997 123 -4951 135
rect -4997 -53 -4991 123
rect -4957 -53 -4951 123
rect -4997 -65 -4951 -53
rect -3339 123 -3293 135
rect -3339 -53 -3333 123
rect -3299 -53 -3293 123
rect -3339 -65 -3293 -53
rect -1681 123 -1635 135
rect -1681 -53 -1675 123
rect -1641 -53 -1635 123
rect -1681 -65 -1635 -53
rect -23 123 23 135
rect -23 -53 -17 123
rect 17 -53 23 123
rect -23 -65 23 -53
rect 1635 123 1681 135
rect 1635 -53 1641 123
rect 1675 -53 1681 123
rect 1635 -65 1681 -53
rect 3293 123 3339 135
rect 3293 -53 3299 123
rect 3333 -53 3339 123
rect 3293 -65 3339 -53
rect 4951 123 4997 135
rect 4951 -53 4957 123
rect 4991 -53 4997 123
rect 4951 -65 4997 -53
rect -4941 -112 -3349 -106
rect -4941 -146 -4929 -112
rect -3361 -146 -3349 -112
rect -4941 -152 -3349 -146
rect -3283 -112 -1691 -106
rect -3283 -146 -3271 -112
rect -1703 -146 -1691 -112
rect -3283 -152 -1691 -146
rect -1625 -112 -33 -106
rect -1625 -146 -1613 -112
rect -45 -146 -33 -112
rect -1625 -152 -33 -146
rect 33 -112 1625 -106
rect 33 -146 45 -112
rect 1613 -146 1625 -112
rect 33 -152 1625 -146
rect 1691 -112 3283 -106
rect 1691 -146 1703 -112
rect 3271 -146 3283 -112
rect 1691 -152 3283 -146
rect 3349 -112 4941 -106
rect 3349 -146 3361 -112
rect 4929 -146 4941 -112
rect 3349 -152 4941 -146
rect -4997 -242 -4951 -230
rect -4997 -418 -4991 -242
rect -4957 -418 -4951 -242
rect -4997 -430 -4951 -418
rect -3339 -242 -3293 -230
rect -3339 -418 -3333 -242
rect -3299 -418 -3293 -242
rect -3339 -430 -3293 -418
rect -1681 -242 -1635 -230
rect -1681 -418 -1675 -242
rect -1641 -418 -1635 -242
rect -1681 -430 -1635 -418
rect -23 -242 23 -230
rect -23 -418 -17 -242
rect 17 -418 23 -242
rect -23 -430 23 -418
rect 1635 -242 1681 -230
rect 1635 -418 1641 -242
rect 1675 -418 1681 -242
rect 1635 -430 1681 -418
rect 3293 -242 3339 -230
rect 3293 -418 3299 -242
rect 3333 -418 3339 -242
rect 3293 -430 3339 -418
rect 4951 -242 4997 -230
rect 4951 -418 4957 -242
rect 4991 -418 4997 -242
rect 4951 -430 4997 -418
rect -4941 -477 -3349 -471
rect -4941 -511 -4929 -477
rect -3361 -511 -3349 -477
rect -4941 -517 -3349 -511
rect -3283 -477 -1691 -471
rect -3283 -511 -3271 -477
rect -1703 -511 -1691 -477
rect -3283 -517 -1691 -511
rect -1625 -477 -33 -471
rect -1625 -511 -1613 -477
rect -45 -511 -33 -477
rect -1625 -517 -33 -511
rect 33 -477 1625 -471
rect 33 -511 45 -477
rect 1613 -511 1625 -477
rect 33 -517 1625 -511
rect 1691 -477 3283 -471
rect 1691 -511 1703 -477
rect 3271 -511 3283 -477
rect 1691 -517 3283 -511
rect 3349 -477 4941 -471
rect 3349 -511 3361 -477
rect 4929 -511 4941 -477
rect 3349 -517 4941 -511
rect -4997 -607 -4951 -595
rect -4997 -783 -4991 -607
rect -4957 -783 -4951 -607
rect -4997 -795 -4951 -783
rect -3339 -607 -3293 -595
rect -3339 -783 -3333 -607
rect -3299 -783 -3293 -607
rect -3339 -795 -3293 -783
rect -1681 -607 -1635 -595
rect -1681 -783 -1675 -607
rect -1641 -783 -1635 -607
rect -1681 -795 -1635 -783
rect -23 -607 23 -595
rect -23 -783 -17 -607
rect 17 -783 23 -607
rect -23 -795 23 -783
rect 1635 -607 1681 -595
rect 1635 -783 1641 -607
rect 1675 -783 1681 -607
rect 1635 -795 1681 -783
rect 3293 -607 3339 -595
rect 3293 -783 3299 -607
rect 3333 -783 3339 -607
rect 3293 -795 3339 -783
rect 4951 -607 4997 -595
rect 4951 -783 4957 -607
rect 4991 -783 4997 -607
rect 4951 -795 4997 -783
rect -4941 -842 -3349 -836
rect -4941 -876 -4929 -842
rect -3361 -876 -3349 -842
rect -4941 -882 -3349 -876
rect -3283 -842 -1691 -836
rect -3283 -876 -3271 -842
rect -1703 -876 -1691 -842
rect -3283 -882 -1691 -876
rect -1625 -842 -33 -836
rect -1625 -876 -1613 -842
rect -45 -876 -33 -842
rect -1625 -882 -33 -876
rect 33 -842 1625 -836
rect 33 -876 45 -842
rect 1613 -876 1625 -842
rect 33 -882 1625 -876
rect 1691 -842 3283 -836
rect 1691 -876 1703 -842
rect 3271 -876 3283 -842
rect 1691 -882 3283 -876
rect 3349 -842 4941 -836
rect 3349 -876 3361 -842
rect 4929 -876 4941 -842
rect 3349 -882 4941 -876
rect -4997 -972 -4951 -960
rect -4997 -1148 -4991 -972
rect -4957 -1148 -4951 -972
rect -4997 -1160 -4951 -1148
rect -3339 -972 -3293 -960
rect -3339 -1148 -3333 -972
rect -3299 -1148 -3293 -972
rect -3339 -1160 -3293 -1148
rect -1681 -972 -1635 -960
rect -1681 -1148 -1675 -972
rect -1641 -1148 -1635 -972
rect -1681 -1160 -1635 -1148
rect -23 -972 23 -960
rect -23 -1148 -17 -972
rect 17 -1148 23 -972
rect -23 -1160 23 -1148
rect 1635 -972 1681 -960
rect 1635 -1148 1641 -972
rect 1675 -1148 1681 -972
rect 1635 -1160 1681 -1148
rect 3293 -972 3339 -960
rect 3293 -1148 3299 -972
rect 3333 -1148 3339 -972
rect 3293 -1160 3339 -1148
rect 4951 -972 4997 -960
rect 4951 -1148 4957 -972
rect 4991 -1148 4997 -972
rect 4951 -1160 4997 -1148
rect -4941 -1207 -3349 -1201
rect -4941 -1241 -4929 -1207
rect -3361 -1241 -3349 -1207
rect -4941 -1247 -3349 -1241
rect -3283 -1207 -1691 -1201
rect -3283 -1241 -3271 -1207
rect -1703 -1241 -1691 -1207
rect -3283 -1247 -1691 -1241
rect -1625 -1207 -33 -1201
rect -1625 -1241 -1613 -1207
rect -45 -1241 -33 -1207
rect -1625 -1247 -33 -1241
rect 33 -1207 1625 -1201
rect 33 -1241 45 -1207
rect 1613 -1241 1625 -1207
rect 33 -1247 1625 -1241
rect 1691 -1207 3283 -1201
rect 1691 -1241 1703 -1207
rect 3271 -1241 3283 -1207
rect 1691 -1247 3283 -1241
rect 3349 -1207 4941 -1201
rect 3349 -1241 3361 -1207
rect 4929 -1241 4941 -1207
rect 3349 -1247 4941 -1241
<< properties >>
string FIXED_BBOX -5108 -1362 5108 1362
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 8 m 7 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712709231
<< pwell >>
rect -2386 -9332 2386 9332
<< psubdiff >>
rect -2350 9262 -2254 9296
rect 2254 9262 2350 9296
rect -2350 9200 -2316 9262
rect 2316 9200 2350 9262
rect -2350 -9262 -2316 -9200
rect 2316 -9262 2350 -9200
rect -2350 -9296 -2254 -9262
rect 2254 -9296 2350 -9262
<< psubdiffcont >>
rect -2254 9262 2254 9296
rect -2350 -9200 -2316 9200
rect 2316 -9200 2350 9200
rect -2254 -9296 2254 -9262
<< xpolycontact >>
rect -2220 8734 -1938 9166
rect -2220 -9166 -1938 -8734
rect -1842 8734 -1560 9166
rect -1842 -9166 -1560 -8734
rect -1464 8734 -1182 9166
rect -1464 -9166 -1182 -8734
rect -1086 8734 -804 9166
rect -1086 -9166 -804 -8734
rect -708 8734 -426 9166
rect -708 -9166 -426 -8734
rect -330 8734 -48 9166
rect -330 -9166 -48 -8734
rect 48 8734 330 9166
rect 48 -9166 330 -8734
rect 426 8734 708 9166
rect 426 -9166 708 -8734
rect 804 8734 1086 9166
rect 804 -9166 1086 -8734
rect 1182 8734 1464 9166
rect 1182 -9166 1464 -8734
rect 1560 8734 1842 9166
rect 1560 -9166 1842 -8734
rect 1938 8734 2220 9166
rect 1938 -9166 2220 -8734
<< xpolyres >>
rect -2220 -8734 -1938 8734
rect -1842 -8734 -1560 8734
rect -1464 -8734 -1182 8734
rect -1086 -8734 -804 8734
rect -708 -8734 -426 8734
rect -330 -8734 -48 8734
rect 48 -8734 330 8734
rect 426 -8734 708 8734
rect 804 -8734 1086 8734
rect 1182 -8734 1464 8734
rect 1560 -8734 1842 8734
rect 1938 -8734 2220 8734
<< locali >>
rect -2350 9262 -2254 9296
rect 2254 9262 2350 9296
rect -2350 9200 -2316 9262
rect 2316 9200 2350 9262
rect -2350 -9262 -2316 -9200
rect 2316 -9262 2350 -9200
rect -2350 -9296 -2254 -9262
rect 2254 -9296 2350 -9262
<< viali >>
rect -2204 8751 -1954 9148
rect -1826 8751 -1576 9148
rect -1448 8751 -1198 9148
rect -1070 8751 -820 9148
rect -692 8751 -442 9148
rect -314 8751 -64 9148
rect 64 8751 314 9148
rect 442 8751 692 9148
rect 820 8751 1070 9148
rect 1198 8751 1448 9148
rect 1576 8751 1826 9148
rect 1954 8751 2204 9148
rect -2204 -9148 -1954 -8751
rect -1826 -9148 -1576 -8751
rect -1448 -9148 -1198 -8751
rect -1070 -9148 -820 -8751
rect -692 -9148 -442 -8751
rect -314 -9148 -64 -8751
rect 64 -9148 314 -8751
rect 442 -9148 692 -8751
rect 820 -9148 1070 -8751
rect 1198 -9148 1448 -8751
rect 1576 -9148 1826 -8751
rect 1954 -9148 2204 -8751
<< metal1 >>
rect -2210 9148 -1948 9160
rect -2210 8751 -2204 9148
rect -1954 8751 -1948 9148
rect -2210 8739 -1948 8751
rect -1832 9148 -1570 9160
rect -1832 8751 -1826 9148
rect -1576 8751 -1570 9148
rect -1832 8739 -1570 8751
rect -1454 9148 -1192 9160
rect -1454 8751 -1448 9148
rect -1198 8751 -1192 9148
rect -1454 8739 -1192 8751
rect -1076 9148 -814 9160
rect -1076 8751 -1070 9148
rect -820 8751 -814 9148
rect -1076 8739 -814 8751
rect -698 9148 -436 9160
rect -698 8751 -692 9148
rect -442 8751 -436 9148
rect -698 8739 -436 8751
rect -320 9148 -58 9160
rect -320 8751 -314 9148
rect -64 8751 -58 9148
rect -320 8739 -58 8751
rect 58 9148 320 9160
rect 58 8751 64 9148
rect 314 8751 320 9148
rect 58 8739 320 8751
rect 436 9148 698 9160
rect 436 8751 442 9148
rect 692 8751 698 9148
rect 436 8739 698 8751
rect 814 9148 1076 9160
rect 814 8751 820 9148
rect 1070 8751 1076 9148
rect 814 8739 1076 8751
rect 1192 9148 1454 9160
rect 1192 8751 1198 9148
rect 1448 8751 1454 9148
rect 1192 8739 1454 8751
rect 1570 9148 1832 9160
rect 1570 8751 1576 9148
rect 1826 8751 1832 9148
rect 1570 8739 1832 8751
rect 1948 9148 2210 9160
rect 1948 8751 1954 9148
rect 2204 8751 2210 9148
rect 1948 8739 2210 8751
rect -2210 -8751 -1948 -8739
rect -2210 -9148 -2204 -8751
rect -1954 -9148 -1948 -8751
rect -2210 -9160 -1948 -9148
rect -1832 -8751 -1570 -8739
rect -1832 -9148 -1826 -8751
rect -1576 -9148 -1570 -8751
rect -1832 -9160 -1570 -9148
rect -1454 -8751 -1192 -8739
rect -1454 -9148 -1448 -8751
rect -1198 -9148 -1192 -8751
rect -1454 -9160 -1192 -9148
rect -1076 -8751 -814 -8739
rect -1076 -9148 -1070 -8751
rect -820 -9148 -814 -8751
rect -1076 -9160 -814 -9148
rect -698 -8751 -436 -8739
rect -698 -9148 -692 -8751
rect -442 -9148 -436 -8751
rect -698 -9160 -436 -9148
rect -320 -8751 -58 -8739
rect -320 -9148 -314 -8751
rect -64 -9148 -58 -8751
rect -320 -9160 -58 -9148
rect 58 -8751 320 -8739
rect 58 -9148 64 -8751
rect 314 -9148 320 -8751
rect 58 -9160 320 -9148
rect 436 -8751 698 -8739
rect 436 -9148 442 -8751
rect 692 -9148 698 -8751
rect 436 -9160 698 -9148
rect 814 -8751 1076 -8739
rect 814 -9148 820 -8751
rect 1070 -9148 1076 -8751
rect 814 -9160 1076 -9148
rect 1192 -8751 1454 -8739
rect 1192 -9148 1198 -8751
rect 1448 -9148 1454 -8751
rect 1192 -9160 1454 -9148
rect 1570 -8751 1832 -8739
rect 1570 -9148 1576 -8751
rect 1826 -9148 1832 -8751
rect 1570 -9160 1832 -9148
rect 1948 -8751 2210 -8739
rect 1948 -9148 1954 -8751
rect 2204 -9148 2210 -8751
rect 1948 -9160 2210 -9148
<< properties >>
string FIXED_BBOX -2333 -9279 2333 9279
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 87.5 m 1 nx 12 wmin 1.410 lmin 0.50 rho 2000 val 124.38k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

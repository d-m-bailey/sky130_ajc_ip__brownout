magic
tech sky130A
magscale 1 2
timestamp 1712352531
<< nwell >>
rect -1374 -797 1374 797
<< mvpmos >>
rect -1116 -500 -716 500
rect -658 -500 -258 500
rect -200 -500 200 500
rect 258 -500 658 500
rect 716 -500 1116 500
<< mvpdiff >>
rect -1174 488 -1116 500
rect -1174 -488 -1162 488
rect -1128 -488 -1116 488
rect -1174 -500 -1116 -488
rect -716 488 -658 500
rect -716 -488 -704 488
rect -670 -488 -658 488
rect -716 -500 -658 -488
rect -258 488 -200 500
rect -258 -488 -246 488
rect -212 -488 -200 488
rect -258 -500 -200 -488
rect 200 488 258 500
rect 200 -488 212 488
rect 246 -488 258 488
rect 200 -500 258 -488
rect 658 488 716 500
rect 658 -488 670 488
rect 704 -488 716 488
rect 658 -500 716 -488
rect 1116 488 1174 500
rect 1116 -488 1128 488
rect 1162 -488 1174 488
rect 1116 -500 1174 -488
<< mvpdiffc >>
rect -1162 -488 -1128 488
rect -704 -488 -670 488
rect -246 -488 -212 488
rect 212 -488 246 488
rect 670 -488 704 488
rect 1128 -488 1162 488
<< mvnsubdiff >>
rect -1308 719 1308 731
rect -1308 685 -1200 719
rect 1200 685 1308 719
rect -1308 673 1308 685
rect -1308 623 -1250 673
rect -1308 -623 -1296 623
rect -1262 -623 -1250 623
rect 1250 623 1308 673
rect -1308 -673 -1250 -623
rect 1250 -623 1262 623
rect 1296 -623 1308 623
rect 1250 -673 1308 -623
rect -1308 -685 1308 -673
rect -1308 -719 -1200 -685
rect 1200 -719 1308 -685
rect -1308 -731 1308 -719
<< mvnsubdiffcont >>
rect -1200 685 1200 719
rect -1296 -623 -1262 623
rect 1262 -623 1296 623
rect -1200 -719 1200 -685
<< poly >>
rect -1116 581 -716 597
rect -1116 547 -1100 581
rect -732 547 -716 581
rect -1116 500 -716 547
rect -658 581 -258 597
rect -658 547 -642 581
rect -274 547 -258 581
rect -658 500 -258 547
rect -200 581 200 597
rect -200 547 -184 581
rect 184 547 200 581
rect -200 500 200 547
rect 258 581 658 597
rect 258 547 274 581
rect 642 547 658 581
rect 258 500 658 547
rect 716 581 1116 597
rect 716 547 732 581
rect 1100 547 1116 581
rect 716 500 1116 547
rect -1116 -547 -716 -500
rect -1116 -581 -1100 -547
rect -732 -581 -716 -547
rect -1116 -597 -716 -581
rect -658 -547 -258 -500
rect -658 -581 -642 -547
rect -274 -581 -258 -547
rect -658 -597 -258 -581
rect -200 -547 200 -500
rect -200 -581 -184 -547
rect 184 -581 200 -547
rect -200 -597 200 -581
rect 258 -547 658 -500
rect 258 -581 274 -547
rect 642 -581 658 -547
rect 258 -597 658 -581
rect 716 -547 1116 -500
rect 716 -581 732 -547
rect 1100 -581 1116 -547
rect 716 -597 1116 -581
<< polycont >>
rect -1100 547 -732 581
rect -642 547 -274 581
rect -184 547 184 581
rect 274 547 642 581
rect 732 547 1100 581
rect -1100 -581 -732 -547
rect -642 -581 -274 -547
rect -184 -581 184 -547
rect 274 -581 642 -547
rect 732 -581 1100 -547
<< locali >>
rect -1296 685 -1200 719
rect 1200 685 1296 719
rect -1296 623 -1262 685
rect 1262 623 1296 685
rect -1116 547 -1100 581
rect -732 547 -716 581
rect -658 547 -642 581
rect -274 547 -258 581
rect -200 547 -184 581
rect 184 547 200 581
rect 258 547 274 581
rect 642 547 658 581
rect 716 547 732 581
rect 1100 547 1116 581
rect -1162 488 -1128 504
rect -1162 -504 -1128 -488
rect -704 488 -670 504
rect -704 -504 -670 -488
rect -246 488 -212 504
rect -246 -504 -212 -488
rect 212 488 246 504
rect 212 -504 246 -488
rect 670 488 704 504
rect 670 -504 704 -488
rect 1128 488 1162 504
rect 1128 -504 1162 -488
rect -1116 -581 -1100 -547
rect -732 -581 -716 -547
rect -658 -581 -642 -547
rect -274 -581 -258 -547
rect -200 -581 -184 -547
rect 184 -581 200 -547
rect 258 -581 274 -547
rect 642 -581 658 -547
rect 716 -581 732 -547
rect 1100 -581 1116 -547
rect -1296 -685 -1262 -623
rect 1262 -685 1296 -623
rect -1296 -719 -1200 -685
rect 1200 -719 1296 -685
<< viali >>
rect -1100 547 -732 581
rect -642 547 -274 581
rect -184 547 184 581
rect 274 547 642 581
rect 732 547 1100 581
rect -1162 -488 -1128 488
rect -704 -488 -670 488
rect -246 -488 -212 488
rect 212 -488 246 488
rect 670 -488 704 488
rect 1128 -488 1162 488
rect -1100 -581 -732 -547
rect -642 -581 -274 -547
rect -184 -581 184 -547
rect 274 -581 642 -547
rect 732 -581 1100 -547
<< metal1 >>
rect -1112 581 -720 587
rect -1112 547 -1100 581
rect -732 547 -720 581
rect -1112 541 -720 547
rect -654 581 -262 587
rect -654 547 -642 581
rect -274 547 -262 581
rect -654 541 -262 547
rect -196 581 196 587
rect -196 547 -184 581
rect 184 547 196 581
rect -196 541 196 547
rect 262 581 654 587
rect 262 547 274 581
rect 642 547 654 581
rect 262 541 654 547
rect 720 581 1112 587
rect 720 547 732 581
rect 1100 547 1112 581
rect 720 541 1112 547
rect -1168 488 -1122 500
rect -1168 -488 -1162 488
rect -1128 -488 -1122 488
rect -1168 -500 -1122 -488
rect -710 488 -664 500
rect -710 -488 -704 488
rect -670 -488 -664 488
rect -710 -500 -664 -488
rect -252 488 -206 500
rect -252 -488 -246 488
rect -212 -488 -206 488
rect -252 -500 -206 -488
rect 206 488 252 500
rect 206 -488 212 488
rect 246 -488 252 488
rect 206 -500 252 -488
rect 664 488 710 500
rect 664 -488 670 488
rect 704 -488 710 488
rect 664 -500 710 -488
rect 1122 488 1168 500
rect 1122 -488 1128 488
rect 1162 -488 1168 488
rect 1122 -500 1168 -488
rect -1112 -547 -720 -541
rect -1112 -581 -1100 -547
rect -732 -581 -720 -547
rect -1112 -587 -720 -581
rect -654 -547 -262 -541
rect -654 -581 -642 -547
rect -274 -581 -262 -547
rect -654 -587 -262 -581
rect -196 -547 196 -541
rect -196 -581 -184 -547
rect 184 -581 196 -547
rect -196 -587 196 -581
rect 262 -547 654 -541
rect 262 -581 274 -547
rect 642 -581 654 -547
rect 262 -587 654 -581
rect 720 -547 1112 -541
rect 720 -581 732 -547
rect 1100 -581 1112 -547
rect 720 -587 1112 -581
<< properties >>
string FIXED_BBOX -1279 -702 1279 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 2 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

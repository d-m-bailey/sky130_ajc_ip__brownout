magic
tech sky130A
magscale 1 2
timestamp 1712554100
<< nwell >>
rect -5203 -677 5203 677
<< mvpmos >>
rect -4945 367 -3345 451
rect -3287 367 -1687 451
rect -1629 367 -29 451
rect 29 367 1629 451
rect 1687 367 3287 451
rect 3345 367 4945 451
rect -4945 118 -3345 202
rect -3287 118 -1687 202
rect -1629 118 -29 202
rect 29 118 1629 202
rect 1687 118 3287 202
rect 3345 118 4945 202
rect -4945 -131 -3345 -47
rect -3287 -131 -1687 -47
rect -1629 -131 -29 -47
rect 29 -131 1629 -47
rect 1687 -131 3287 -47
rect 3345 -131 4945 -47
rect -4945 -380 -3345 -296
rect -3287 -380 -1687 -296
rect -1629 -380 -29 -296
rect 29 -380 1629 -296
rect 1687 -380 3287 -296
rect 3345 -380 4945 -296
<< mvpdiff >>
rect -5003 439 -4945 451
rect -5003 379 -4991 439
rect -4957 379 -4945 439
rect -5003 367 -4945 379
rect -3345 439 -3287 451
rect -3345 379 -3333 439
rect -3299 379 -3287 439
rect -3345 367 -3287 379
rect -1687 439 -1629 451
rect -1687 379 -1675 439
rect -1641 379 -1629 439
rect -1687 367 -1629 379
rect -29 439 29 451
rect -29 379 -17 439
rect 17 379 29 439
rect -29 367 29 379
rect 1629 439 1687 451
rect 1629 379 1641 439
rect 1675 379 1687 439
rect 1629 367 1687 379
rect 3287 439 3345 451
rect 3287 379 3299 439
rect 3333 379 3345 439
rect 3287 367 3345 379
rect 4945 439 5003 451
rect 4945 379 4957 439
rect 4991 379 5003 439
rect 4945 367 5003 379
rect -5003 190 -4945 202
rect -5003 130 -4991 190
rect -4957 130 -4945 190
rect -5003 118 -4945 130
rect -3345 190 -3287 202
rect -3345 130 -3333 190
rect -3299 130 -3287 190
rect -3345 118 -3287 130
rect -1687 190 -1629 202
rect -1687 130 -1675 190
rect -1641 130 -1629 190
rect -1687 118 -1629 130
rect -29 190 29 202
rect -29 130 -17 190
rect 17 130 29 190
rect -29 118 29 130
rect 1629 190 1687 202
rect 1629 130 1641 190
rect 1675 130 1687 190
rect 1629 118 1687 130
rect 3287 190 3345 202
rect 3287 130 3299 190
rect 3333 130 3345 190
rect 3287 118 3345 130
rect 4945 190 5003 202
rect 4945 130 4957 190
rect 4991 130 5003 190
rect 4945 118 5003 130
rect -5003 -59 -4945 -47
rect -5003 -119 -4991 -59
rect -4957 -119 -4945 -59
rect -5003 -131 -4945 -119
rect -3345 -59 -3287 -47
rect -3345 -119 -3333 -59
rect -3299 -119 -3287 -59
rect -3345 -131 -3287 -119
rect -1687 -59 -1629 -47
rect -1687 -119 -1675 -59
rect -1641 -119 -1629 -59
rect -1687 -131 -1629 -119
rect -29 -59 29 -47
rect -29 -119 -17 -59
rect 17 -119 29 -59
rect -29 -131 29 -119
rect 1629 -59 1687 -47
rect 1629 -119 1641 -59
rect 1675 -119 1687 -59
rect 1629 -131 1687 -119
rect 3287 -59 3345 -47
rect 3287 -119 3299 -59
rect 3333 -119 3345 -59
rect 3287 -131 3345 -119
rect 4945 -59 5003 -47
rect 4945 -119 4957 -59
rect 4991 -119 5003 -59
rect 4945 -131 5003 -119
rect -5003 -308 -4945 -296
rect -5003 -368 -4991 -308
rect -4957 -368 -4945 -308
rect -5003 -380 -4945 -368
rect -3345 -308 -3287 -296
rect -3345 -368 -3333 -308
rect -3299 -368 -3287 -308
rect -3345 -380 -3287 -368
rect -1687 -308 -1629 -296
rect -1687 -368 -1675 -308
rect -1641 -368 -1629 -308
rect -1687 -380 -1629 -368
rect -29 -308 29 -296
rect -29 -368 -17 -308
rect 17 -368 29 -308
rect -29 -380 29 -368
rect 1629 -308 1687 -296
rect 1629 -368 1641 -308
rect 1675 -368 1687 -308
rect 1629 -380 1687 -368
rect 3287 -308 3345 -296
rect 3287 -368 3299 -308
rect 3333 -368 3345 -308
rect 3287 -380 3345 -368
rect 4945 -308 5003 -296
rect 4945 -368 4957 -308
rect 4991 -368 5003 -308
rect 4945 -380 5003 -368
<< mvpdiffc >>
rect -4991 379 -4957 439
rect -3333 379 -3299 439
rect -1675 379 -1641 439
rect -17 379 17 439
rect 1641 379 1675 439
rect 3299 379 3333 439
rect 4957 379 4991 439
rect -4991 130 -4957 190
rect -3333 130 -3299 190
rect -1675 130 -1641 190
rect -17 130 17 190
rect 1641 130 1675 190
rect 3299 130 3333 190
rect 4957 130 4991 190
rect -4991 -119 -4957 -59
rect -3333 -119 -3299 -59
rect -1675 -119 -1641 -59
rect -17 -119 17 -59
rect 1641 -119 1675 -59
rect 3299 -119 3333 -59
rect 4957 -119 4991 -59
rect -4991 -368 -4957 -308
rect -3333 -368 -3299 -308
rect -1675 -368 -1641 -308
rect -17 -368 17 -308
rect 1641 -368 1675 -308
rect 3299 -368 3333 -308
rect 4957 -368 4991 -308
<< mvnsubdiff >>
rect -5137 599 5137 611
rect -5137 565 -5029 599
rect 5029 565 5137 599
rect -5137 553 5137 565
rect -5137 503 -5079 553
rect -5137 -503 -5125 503
rect -5091 -503 -5079 503
rect 5079 503 5137 553
rect -5137 -553 -5079 -503
rect 5079 -503 5091 503
rect 5125 -503 5137 503
rect 5079 -553 5137 -503
rect -5137 -565 5137 -553
rect -5137 -599 -5029 -565
rect 5029 -599 5137 -565
rect -5137 -611 5137 -599
<< mvnsubdiffcont >>
rect -5029 565 5029 599
rect -5125 -503 -5091 503
rect 5091 -503 5125 503
rect -5029 -599 5029 -565
<< poly >>
rect -4945 451 -3345 477
rect -3287 451 -1687 477
rect -1629 451 -29 477
rect 29 451 1629 477
rect 1687 451 3287 477
rect 3345 451 4945 477
rect -4945 320 -3345 367
rect -4945 286 -4929 320
rect -3361 286 -3345 320
rect -4945 270 -3345 286
rect -3287 320 -1687 367
rect -3287 286 -3271 320
rect -1703 286 -1687 320
rect -3287 270 -1687 286
rect -1629 320 -29 367
rect -1629 286 -1613 320
rect -45 286 -29 320
rect -1629 270 -29 286
rect 29 320 1629 367
rect 29 286 45 320
rect 1613 286 1629 320
rect 29 270 1629 286
rect 1687 320 3287 367
rect 1687 286 1703 320
rect 3271 286 3287 320
rect 1687 270 3287 286
rect 3345 320 4945 367
rect 3345 286 3361 320
rect 4929 286 4945 320
rect 3345 270 4945 286
rect -4945 202 -3345 228
rect -3287 202 -1687 228
rect -1629 202 -29 228
rect 29 202 1629 228
rect 1687 202 3287 228
rect 3345 202 4945 228
rect -4945 71 -3345 118
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -4945 21 -3345 37
rect -3287 71 -1687 118
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -3287 21 -1687 37
rect -1629 71 -29 118
rect -1629 37 -1613 71
rect -45 37 -29 71
rect -1629 21 -29 37
rect 29 71 1629 118
rect 29 37 45 71
rect 1613 37 1629 71
rect 29 21 1629 37
rect 1687 71 3287 118
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 1687 21 3287 37
rect 3345 71 4945 118
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 3345 21 4945 37
rect -4945 -47 -3345 -21
rect -3287 -47 -1687 -21
rect -1629 -47 -29 -21
rect 29 -47 1629 -21
rect 1687 -47 3287 -21
rect 3345 -47 4945 -21
rect -4945 -178 -3345 -131
rect -4945 -212 -4929 -178
rect -3361 -212 -3345 -178
rect -4945 -228 -3345 -212
rect -3287 -178 -1687 -131
rect -3287 -212 -3271 -178
rect -1703 -212 -1687 -178
rect -3287 -228 -1687 -212
rect -1629 -178 -29 -131
rect -1629 -212 -1613 -178
rect -45 -212 -29 -178
rect -1629 -228 -29 -212
rect 29 -178 1629 -131
rect 29 -212 45 -178
rect 1613 -212 1629 -178
rect 29 -228 1629 -212
rect 1687 -178 3287 -131
rect 1687 -212 1703 -178
rect 3271 -212 3287 -178
rect 1687 -228 3287 -212
rect 3345 -178 4945 -131
rect 3345 -212 3361 -178
rect 4929 -212 4945 -178
rect 3345 -228 4945 -212
rect -4945 -296 -3345 -270
rect -3287 -296 -1687 -270
rect -1629 -296 -29 -270
rect 29 -296 1629 -270
rect 1687 -296 3287 -270
rect 3345 -296 4945 -270
rect -4945 -427 -3345 -380
rect -4945 -461 -4929 -427
rect -3361 -461 -3345 -427
rect -4945 -477 -3345 -461
rect -3287 -427 -1687 -380
rect -3287 -461 -3271 -427
rect -1703 -461 -1687 -427
rect -3287 -477 -1687 -461
rect -1629 -427 -29 -380
rect -1629 -461 -1613 -427
rect -45 -461 -29 -427
rect -1629 -477 -29 -461
rect 29 -427 1629 -380
rect 29 -461 45 -427
rect 1613 -461 1629 -427
rect 29 -477 1629 -461
rect 1687 -427 3287 -380
rect 1687 -461 1703 -427
rect 3271 -461 3287 -427
rect 1687 -477 3287 -461
rect 3345 -427 4945 -380
rect 3345 -461 3361 -427
rect 4929 -461 4945 -427
rect 3345 -477 4945 -461
<< polycont >>
rect -4929 286 -3361 320
rect -3271 286 -1703 320
rect -1613 286 -45 320
rect 45 286 1613 320
rect 1703 286 3271 320
rect 3361 286 4929 320
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect -4929 -212 -3361 -178
rect -3271 -212 -1703 -178
rect -1613 -212 -45 -178
rect 45 -212 1613 -178
rect 1703 -212 3271 -178
rect 3361 -212 4929 -178
rect -4929 -461 -3361 -427
rect -3271 -461 -1703 -427
rect -1613 -461 -45 -427
rect 45 -461 1613 -427
rect 1703 -461 3271 -427
rect 3361 -461 4929 -427
<< locali >>
rect -5125 565 -5029 599
rect 5029 565 5125 599
rect -5125 503 -5091 565
rect 5091 503 5125 565
rect -4991 439 -4957 455
rect -4991 363 -4957 379
rect -3333 439 -3299 455
rect -3333 363 -3299 379
rect -1675 439 -1641 455
rect -1675 363 -1641 379
rect -17 439 17 455
rect -17 363 17 379
rect 1641 439 1675 455
rect 1641 363 1675 379
rect 3299 439 3333 455
rect 3299 363 3333 379
rect 4957 439 4991 455
rect 4957 363 4991 379
rect -4945 286 -4929 320
rect -3361 286 -3345 320
rect -3287 286 -3271 320
rect -1703 286 -1687 320
rect -1629 286 -1613 320
rect -45 286 -29 320
rect 29 286 45 320
rect 1613 286 1629 320
rect 1687 286 1703 320
rect 3271 286 3287 320
rect 3345 286 3361 320
rect 4929 286 4945 320
rect -4991 190 -4957 206
rect -4991 114 -4957 130
rect -3333 190 -3299 206
rect -3333 114 -3299 130
rect -1675 190 -1641 206
rect -1675 114 -1641 130
rect -17 190 17 206
rect -17 114 17 130
rect 1641 190 1675 206
rect 1641 114 1675 130
rect 3299 190 3333 206
rect 3299 114 3333 130
rect 4957 190 4991 206
rect 4957 114 4991 130
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -1629 37 -1613 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1613 37 1629 71
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 3345 37 3361 71
rect 4929 37 4945 71
rect -4991 -59 -4957 -43
rect -4991 -135 -4957 -119
rect -3333 -59 -3299 -43
rect -3333 -135 -3299 -119
rect -1675 -59 -1641 -43
rect -1675 -135 -1641 -119
rect -17 -59 17 -43
rect -17 -135 17 -119
rect 1641 -59 1675 -43
rect 1641 -135 1675 -119
rect 3299 -59 3333 -43
rect 3299 -135 3333 -119
rect 4957 -59 4991 -43
rect 4957 -135 4991 -119
rect -4945 -212 -4929 -178
rect -3361 -212 -3345 -178
rect -3287 -212 -3271 -178
rect -1703 -212 -1687 -178
rect -1629 -212 -1613 -178
rect -45 -212 -29 -178
rect 29 -212 45 -178
rect 1613 -212 1629 -178
rect 1687 -212 1703 -178
rect 3271 -212 3287 -178
rect 3345 -212 3361 -178
rect 4929 -212 4945 -178
rect -4991 -308 -4957 -292
rect -4991 -384 -4957 -368
rect -3333 -308 -3299 -292
rect -3333 -384 -3299 -368
rect -1675 -308 -1641 -292
rect -1675 -384 -1641 -368
rect -17 -308 17 -292
rect -17 -384 17 -368
rect 1641 -308 1675 -292
rect 1641 -384 1675 -368
rect 3299 -308 3333 -292
rect 3299 -384 3333 -368
rect 4957 -308 4991 -292
rect 4957 -384 4991 -368
rect -4945 -461 -4929 -427
rect -3361 -461 -3345 -427
rect -3287 -461 -3271 -427
rect -1703 -461 -1687 -427
rect -1629 -461 -1613 -427
rect -45 -461 -29 -427
rect 29 -461 45 -427
rect 1613 -461 1629 -427
rect 1687 -461 1703 -427
rect 3271 -461 3287 -427
rect 3345 -461 3361 -427
rect 4929 -461 4945 -427
rect -5125 -565 -5091 -503
rect 5091 -565 5125 -503
rect -5125 -599 -5029 -565
rect 5029 -599 5125 -565
<< viali >>
rect -4991 379 -4957 439
rect -3333 379 -3299 439
rect -1675 379 -1641 439
rect -17 379 17 439
rect 1641 379 1675 439
rect 3299 379 3333 439
rect 4957 379 4991 439
rect -4929 286 -3361 320
rect -3271 286 -1703 320
rect -1613 286 -45 320
rect 45 286 1613 320
rect 1703 286 3271 320
rect 3361 286 4929 320
rect -4991 130 -4957 190
rect -3333 130 -3299 190
rect -1675 130 -1641 190
rect -17 130 17 190
rect 1641 130 1675 190
rect 3299 130 3333 190
rect 4957 130 4991 190
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect -4991 -119 -4957 -59
rect -3333 -119 -3299 -59
rect -1675 -119 -1641 -59
rect -17 -119 17 -59
rect 1641 -119 1675 -59
rect 3299 -119 3333 -59
rect 4957 -119 4991 -59
rect -4929 -212 -3361 -178
rect -3271 -212 -1703 -178
rect -1613 -212 -45 -178
rect 45 -212 1613 -178
rect 1703 -212 3271 -178
rect 3361 -212 4929 -178
rect -4991 -368 -4957 -308
rect -3333 -368 -3299 -308
rect -1675 -368 -1641 -308
rect -17 -368 17 -308
rect 1641 -368 1675 -308
rect 3299 -368 3333 -308
rect 4957 -368 4991 -308
rect -4929 -461 -3361 -427
rect -3271 -461 -1703 -427
rect -1613 -461 -45 -427
rect 45 -461 1613 -427
rect 1703 -461 3271 -427
rect 3361 -461 4929 -427
<< metal1 >>
rect -4997 439 -4951 451
rect -4997 379 -4991 439
rect -4957 379 -4951 439
rect -4997 367 -4951 379
rect -3339 439 -3293 451
rect -3339 379 -3333 439
rect -3299 379 -3293 439
rect -3339 367 -3293 379
rect -1681 439 -1635 451
rect -1681 379 -1675 439
rect -1641 379 -1635 439
rect -1681 367 -1635 379
rect -23 439 23 451
rect -23 379 -17 439
rect 17 379 23 439
rect -23 367 23 379
rect 1635 439 1681 451
rect 1635 379 1641 439
rect 1675 379 1681 439
rect 1635 367 1681 379
rect 3293 439 3339 451
rect 3293 379 3299 439
rect 3333 379 3339 439
rect 3293 367 3339 379
rect 4951 439 4997 451
rect 4951 379 4957 439
rect 4991 379 4997 439
rect 4951 367 4997 379
rect -4941 320 -3349 326
rect -4941 286 -4929 320
rect -3361 286 -3349 320
rect -4941 280 -3349 286
rect -3283 320 -1691 326
rect -3283 286 -3271 320
rect -1703 286 -1691 320
rect -3283 280 -1691 286
rect -1625 320 -33 326
rect -1625 286 -1613 320
rect -45 286 -33 320
rect -1625 280 -33 286
rect 33 320 1625 326
rect 33 286 45 320
rect 1613 286 1625 320
rect 33 280 1625 286
rect 1691 320 3283 326
rect 1691 286 1703 320
rect 3271 286 3283 320
rect 1691 280 3283 286
rect 3349 320 4941 326
rect 3349 286 3361 320
rect 4929 286 4941 320
rect 3349 280 4941 286
rect -4997 190 -4951 202
rect -4997 130 -4991 190
rect -4957 130 -4951 190
rect -4997 118 -4951 130
rect -3339 190 -3293 202
rect -3339 130 -3333 190
rect -3299 130 -3293 190
rect -3339 118 -3293 130
rect -1681 190 -1635 202
rect -1681 130 -1675 190
rect -1641 130 -1635 190
rect -1681 118 -1635 130
rect -23 190 23 202
rect -23 130 -17 190
rect 17 130 23 190
rect -23 118 23 130
rect 1635 190 1681 202
rect 1635 130 1641 190
rect 1675 130 1681 190
rect 1635 118 1681 130
rect 3293 190 3339 202
rect 3293 130 3299 190
rect 3333 130 3339 190
rect 3293 118 3339 130
rect 4951 190 4997 202
rect 4951 130 4957 190
rect 4991 130 4997 190
rect 4951 118 4997 130
rect -4941 71 -3349 77
rect -4941 37 -4929 71
rect -3361 37 -3349 71
rect -4941 31 -3349 37
rect -3283 71 -1691 77
rect -3283 37 -3271 71
rect -1703 37 -1691 71
rect -3283 31 -1691 37
rect -1625 71 -33 77
rect -1625 37 -1613 71
rect -45 37 -33 71
rect -1625 31 -33 37
rect 33 71 1625 77
rect 33 37 45 71
rect 1613 37 1625 71
rect 33 31 1625 37
rect 1691 71 3283 77
rect 1691 37 1703 71
rect 3271 37 3283 71
rect 1691 31 3283 37
rect 3349 71 4941 77
rect 3349 37 3361 71
rect 4929 37 4941 71
rect 3349 31 4941 37
rect -4997 -59 -4951 -47
rect -4997 -119 -4991 -59
rect -4957 -119 -4951 -59
rect -4997 -131 -4951 -119
rect -3339 -59 -3293 -47
rect -3339 -119 -3333 -59
rect -3299 -119 -3293 -59
rect -3339 -131 -3293 -119
rect -1681 -59 -1635 -47
rect -1681 -119 -1675 -59
rect -1641 -119 -1635 -59
rect -1681 -131 -1635 -119
rect -23 -59 23 -47
rect -23 -119 -17 -59
rect 17 -119 23 -59
rect -23 -131 23 -119
rect 1635 -59 1681 -47
rect 1635 -119 1641 -59
rect 1675 -119 1681 -59
rect 1635 -131 1681 -119
rect 3293 -59 3339 -47
rect 3293 -119 3299 -59
rect 3333 -119 3339 -59
rect 3293 -131 3339 -119
rect 4951 -59 4997 -47
rect 4951 -119 4957 -59
rect 4991 -119 4997 -59
rect 4951 -131 4997 -119
rect -4941 -178 -3349 -172
rect -4941 -212 -4929 -178
rect -3361 -212 -3349 -178
rect -4941 -218 -3349 -212
rect -3283 -178 -1691 -172
rect -3283 -212 -3271 -178
rect -1703 -212 -1691 -178
rect -3283 -218 -1691 -212
rect -1625 -178 -33 -172
rect -1625 -212 -1613 -178
rect -45 -212 -33 -178
rect -1625 -218 -33 -212
rect 33 -178 1625 -172
rect 33 -212 45 -178
rect 1613 -212 1625 -178
rect 33 -218 1625 -212
rect 1691 -178 3283 -172
rect 1691 -212 1703 -178
rect 3271 -212 3283 -178
rect 1691 -218 3283 -212
rect 3349 -178 4941 -172
rect 3349 -212 3361 -178
rect 4929 -212 4941 -178
rect 3349 -218 4941 -212
rect -4997 -308 -4951 -296
rect -4997 -368 -4991 -308
rect -4957 -368 -4951 -308
rect -4997 -380 -4951 -368
rect -3339 -308 -3293 -296
rect -3339 -368 -3333 -308
rect -3299 -368 -3293 -308
rect -3339 -380 -3293 -368
rect -1681 -308 -1635 -296
rect -1681 -368 -1675 -308
rect -1641 -368 -1635 -308
rect -1681 -380 -1635 -368
rect -23 -308 23 -296
rect -23 -368 -17 -308
rect 17 -368 23 -308
rect -23 -380 23 -368
rect 1635 -308 1681 -296
rect 1635 -368 1641 -308
rect 1675 -368 1681 -308
rect 1635 -380 1681 -368
rect 3293 -308 3339 -296
rect 3293 -368 3299 -308
rect 3333 -368 3339 -308
rect 3293 -380 3339 -368
rect 4951 -308 4997 -296
rect 4951 -368 4957 -308
rect 4991 -368 4997 -308
rect 4951 -380 4997 -368
rect -4941 -427 -3349 -421
rect -4941 -461 -4929 -427
rect -3361 -461 -3349 -427
rect -4941 -467 -3349 -461
rect -3283 -427 -1691 -421
rect -3283 -461 -3271 -427
rect -1703 -461 -1691 -427
rect -3283 -467 -1691 -461
rect -1625 -427 -33 -421
rect -1625 -461 -1613 -427
rect -45 -461 -33 -427
rect -1625 -467 -33 -461
rect 33 -427 1625 -421
rect 33 -461 45 -427
rect 1613 -461 1625 -427
rect 33 -467 1625 -461
rect 1691 -427 3283 -421
rect 1691 -461 1703 -427
rect 3271 -461 3283 -427
rect 1691 -467 3283 -461
rect 3349 -427 4941 -421
rect 3349 -461 3361 -427
rect 4929 -461 4941 -427
rect 3349 -467 4941 -461
<< properties >>
string FIXED_BBOX -5108 -582 5108 582
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8 m 4 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

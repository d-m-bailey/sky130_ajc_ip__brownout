* NGSPICE file created from brownout_ana_rcx.ext - technology: sky130A

*.subckt brownout_ana_rcx otrip_decoded[1] otrip_decoded[0] vin_vunder ena ibg_200n
*+ itest vtrip_decoded[6] vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2]
*+ vtrip_decoded[0] osc_ck outb otrip_decoded[7] vunder otrip_decoded[4] isrc_sel otrip_decoded[5]
*+ otrip_decoded[2] vbg_1v2 vin_brout brout_filt dcomp outb_unbuf vtrip_decoded[7]
*+ vtrip_decoded[1] otrip_decoded[3] otrip_decoded[6] avss dvdd dvss avdd osc_ena

.subckt brownout_ana vin_brout otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3]
+ otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vin_vunder vbg_1v2 ena avdd ibg_200n itest avss dvdd isrc_sel dvss vtrip_decoded[7]
+ vtrip_decoded[6] vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2] vtrip_decoded[1] vtrip_decoded[0] dcomp brout_filt osc_ck
+ osc_ena vunder outb outb_unbuf

X0 a_8447_n11914# a_8069_n19314# avss.t101 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 avss.t357 comparator_1.n1 dcomp3v3 avss.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X2 comparator_1.vt avss.t366 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X3 a_n15745_n11914# a_n16123_n19314# avss.t99 sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 rstring_mux_0.vtrip4.t4 rstring_mux_0.vtrip_decoded_avdd[4] vin_vunder.t23 avss.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 avdd.t601 comparator_1.n1 dcomp3v3 avdd.t600 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X6 dvdd.t277 sky130_fd_sc_hd__inv_4_1.Y vunder.t2 dvdd.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 rstring_mux_0.vtrip_decoded_b_avdd[7] rstring_mux_0.vtrip_decoded_avdd[7] avss.t308 avss.t307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X8 dvdd.t126 dvdd.t124 osc_ck.t4 dvdd.t125 sky130_fd_pr__pfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X9 a_5346_n3990# a_4921_n3946# dvss.t651 dvss.t650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X10 rc_osc_0.n.t0 dvdd.t122 rc_osc_0.m dvdd.t123 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 dvdd.t39 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t15 dvdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 avdd.t115 a_429_n2876# a_1122_n3990# avdd.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X13 rstring_mux_0.vtop.t17 a_n16123_n19314# avss.t185 sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 comparator_0.vn comparator_0.ena comparator_0.ibias avss.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X15 avss.t97 avss.t96 avss.t97 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X16 dvss.t51 otrip_decoded[0].t0 a_n8119_n2964# dvss.t50 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X17 comparator_1.vpp comparator_0.ena avdd.t562 avdd.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X18 comparator_1.n0 comparator_1.vpp avdd.t481 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X19 dvss.t354 a_7033_n3946# a_7458_n3990# dvss.t353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X20 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.otrip_decoded_avdd[1] avss.t190 avss.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X21 vin_brout avdd.t400 vin_brout avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=23.2 ps=169.28 w=5 l=0.6
X22 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 comparator_1.vpp comparator_1.vnn avdd.t150 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X24 dcomp.t15 sky130_fd_sc_hd__inv_4_3.Y dvdd.t321 dvdd.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 dvdd.t81 schmitt_trigger_0.in.t1 schmitt_trigger_0.m.t5 dvdd.t80 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 comparator_0.vnn vin_vunder.t48 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X27 a_3155_n11914# a_3533_n19314# avss.t215 sky130_fd_pr__res_xhigh_po_1p41 l=35
X28 a_n11209_n11914# a_n10831_n19314# avss.t167 sky130_fd_pr__res_xhigh_po_1p41 l=35
X29 comparator_1.vpp vbg_1v2.t0 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X30 rstring_mux_0.otrip_decoded_avdd[5] a_n2588_n1478# avdd.t576 avdd.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X31 dvdd.t7 a_10873_n2760# a_10873_n3956# dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X32 a_7458_n3990# a_7033_n3946# dvss.t352 dvss.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X33 comparator_1.vpp comparator_1.vnn avdd.t149 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X34 ibias_gen_0.vr.t3 ibias_gen_0.vn0.t19 ibias_gen_0.vp0.t2 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X35 avdd.t57 a_2541_n2876# a_3234_n3990# avdd.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X36 comparator_0.vpp comparator_0.vnn avdd.t204 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X37 a_n26830_n2937# a_n27208_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X38 dvdd.t166 sky130_fd_sc_hd__inv_4_4.Y outb.t15 dvdd.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X39 dvss.t158 a_9145_n3946# a_9570_n3990# dvss.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X40 comparator_0.vt vin_vunder.t49 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X41 rstring_mux_0.vtrip_decoded_avdd[0] a_1636_n3212# dvss.t597 dvss.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X42 dvss.t15 a_6765_n2876# a_7972_n3212# dvss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X43 avdd.t575 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b avdd.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X44 a_n8951_9395# a_n8573_1995# avss.t100 sky130_fd_pr__res_xhigh_po_1p41 l=35
X45 itest.t1 ibias_gen_0.vp.t7 avdd.t91 avdd.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X46 vin_vunder.t43 avdd.t398 vin_vunder.t43 avdd.t399 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X47 comparator_1.vt vbg_1v2.t1 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X48 rstring_mux_0.vtrip7.t1 a_n247_n19314# avss.t119 sky130_fd_pr__res_xhigh_po_1p41 l=35
X49 dvss.t93 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t31 dvss.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X50 comparator_1.vt vbg_1v2.t2 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X51 a_n24562_n2937# a_n24184_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X52 a_n21538_n2937# a_n21160_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X53 avdd.t608 a_4653_n2876# a_5346_n3990# avdd.t607 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X54 vin_brout avdd.t396 vin_brout avdd.t397 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X55 dvdd.t164 sky130_fd_sc_hd__inv_4_4.Y outb.t14 dvdd.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X56 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.otrip_decoded_avdd[2] avss.t138 avss.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X57 a_6935_n11914# a_6557_n19314# avss.t193 sky130_fd_pr__res_xhigh_po_1p41 l=35
X58 avss.t301 comparator_0.ena rstring_mux_0.ena_b avss.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X59 a_n26830_n2937# a_n26452_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X60 a_n23806_n2937# a_n23428_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X61 comparator_0.vpp comparator_0.vnn avdd.t203 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X62 rstring_mux_0.vtrip2.t9 rstring_mux_0.vtrip_decoded_avdd[2] vin_vunder.t19 avss.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X63 outb.t31 sky130_fd_sc_hd__inv_4_4.Y dvss.t417 dvss.t416 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X64 rstring_mux_0.vtrip_decoded_avdd[2] a_3748_n3212# dvss.t358 dvss.t357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X65 a_n7326_n3990# a_n7751_n3946# dvss.t11 dvss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X66 a_6935_n11914# a_7313_n19314# avss.t116 sky130_fd_pr__res_xhigh_po_1p41 l=35
X67 a_n14989_n11914# a_n14611_n19314# avss.t179 sky130_fd_pr__res_xhigh_po_1p41 l=35
X68 a_n3649_n11914# a_n4027_n19314# avss.t130 sky130_fd_pr__res_xhigh_po_1p41 l=35
X69 dvdd.t73 vl sky130_fd_sc_hd__inv_4_3.Y dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X70 avdd.t455 a_n3795_n1142# a_n2588_n1478# avdd.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X71 dvss.t730 sky130_fd_sc_hd__inv_4_3.Y dcomp.t31 dvss.t729 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 comparator_0.vnn comparator_0.vpp avdd.t45 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X73 a_n4405_n11914# a_n4027_n19314# avss.t178 sky130_fd_pr__res_xhigh_po_1p41 l=35
X74 ibias_gen_0.vp1.t9 ibias_gen_0.vp1.t8 avdd.t449 avdd.t448 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X75 a_n15529_n2223# ibias_gen_0.isrc_sel_b ibias_gen_0.vn1.t7 avdd.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X76 a_n1683_n1142# a_n1783_n1230# dvss.t120 dvss.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X77 dvss.t641 vtrip_decoded[3].t0 a_2441_n1230# dvss.t640 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X78 comparator_0.vpp comparator_0.vnn avdd.t202 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X79 avdd.t210 a_n3102_n2256# a_n3795_n1142# avdd.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X80 avdd.t13 a_6765_n2876# a_7458_n3990# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X81 a_2809_n3946# a_2441_n2964# dvdd.t239 dvdd.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X82 dvdd.t162 sky130_fd_sc_hd__inv_4_4.Y outb.t13 dvdd.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X83 dvdd.t275 sky130_fd_sc_hd__inv_4_1.Y vunder.t8 dvdd.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X84 dvss.t108 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X sky130_fd_sc_hd__inv_4_1.A dvss.t107 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X85 osc_ck.t5 osc_ena.t0 rc_osc_0.vr dvss.t383 sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X86 avdd.t201 comparator_0.vnn comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X87 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.otrip_decoded_avdd[6] avdd.t208 avdd.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X88 a_n10279_n24223# a_11121_n24601# dvss.t523 sky130_fd_pr__res_xhigh_po_1p41 l=105
X89 dcomp.t14 sky130_fd_sc_hd__inv_4_3.Y dvdd.t319 dvdd.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 dvdd.t37 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t14 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X91 rstring_mux_0.vtrip3.t6 rstring_mux_0.vtrip_decoded_b_avdd[3] vin_vunder.t34 avdd.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X92 dvdd.t287 rc_osc_0.m rc_osc_0.n.t3 dvdd.t286 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X93 avss.t286 comparator_1.vn comparator_1.vn avss.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X94 ibias_gen_0.vn0.t15 vbg_1v2.t3 ibias_gen_0.vstart.t10 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X95 rc_osc_0.m rc_osc_0.in dvdd.t194 dvdd.t193 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X96 ibias_gen_0.vr.t4 a_n20404_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X97 avdd.t521 a_n5907_n1142# a_n4700_n1478# avdd.t517 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X98 comparator_1.ena_b comparator_0.ena avdd.t560 avdd.t559 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X99 dvss.t629 sky130_fd_sc_hd__inv_4_1.Y vunder.t31 dvss.t628 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X100 a_n13487_9395# a_n13109_1995# avss.t184 sky130_fd_pr__res_xhigh_po_1p41 l=35
X101 a_n3795_n1142# a_n3895_n1230# dvss.t265 dvss.t264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X102 a_2541_n1142# a_2441_n1230# dvss.t581 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X103 a_7033_n3946# a_6665_n2964# dvdd.t243 dvdd.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X104 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvss.t553 dvss.t552 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X105 schmitt_trigger_0.m.t8 schmitt_trigger_0.out.t4 dvdd.t101 dvdd.t100 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X106 a_n14243_9395# a_n14621_1995# avss.t118 sky130_fd_pr__res_xhigh_po_1p41 l=35
X107 dvdd.t121 dvdd.t119 schmitt_trigger_0.m.t12 dvdd.t120 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X108 dvdd.t5 otrip_decoded[6].t0 a_n1783_n2964# dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X109 avss.t355 comparator_1.n1 dcomp3v3 avss.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X110 dvss.t100 a_8877_n1142# a_10084_n1478# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X111 rstring_mux_0.vtrip_decoded_avdd[5] a_5860_n1478# avdd.t525 avdd.t515 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X112 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.otrip_decoded_avdd[1] avdd.t212 avdd.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X113 a_n7429_n11914# a_n7807_n19314# avss.t122 sky130_fd_pr__res_xhigh_po_1p41 l=35
X114 dvss.t122 a_2541_n2876# a_3748_n3212# dvss.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X115 comparator_0.vnn comparator_0.vpp avdd.t44 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X116 avdd.t161 a_n8019_n1142# a_n6812_n1478# avdd.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X117 dcomp3v3uv comparator_0.n1 avdd.t439 avdd.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X118 vin_vunder.t21 rstring_mux_0.vtrip_decoded_b_avdd[5] rstring_mux_0.vtrip5.t7 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X119 rstring_mux_0.otrip_decoded_avdd[5] a_n2588_n1478# dvss.t697 dvss.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X120 avdd.t480 comparator_1.vpp comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X121 a_4653_n1142# a_4553_n1230# dvss.t533 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X122 a_9145_n3946# a_8777_n2964# dvdd.t128 dvdd.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X123 avdd.t200 comparator_0.vnn comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X124 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X125 a_5423_n11914# a_5801_n19314# avss.t222 sky130_fd_pr__res_xhigh_po_1p41 l=35
X126 avdd.t148 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X127 comparator_0.vnn vin_vunder.t50 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X128 dvss.t448 outb_unbuf.t0 sky130_fd_sc_hd__inv_4_4.Y dvss.t447 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 dvdd.t210 otrip_decoded[4].t0 a_n3895_n2964# dvdd.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X130 a_n11975_9395# a_n11597_1995# avss.t117 sky130_fd_pr__res_xhigh_po_1p41 l=35
X131 dvss.t91 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t30 dvss.t90 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X132 dvss.t97 vtrip_decoded[1].t0 a_329_n1230# dvss.t96 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X133 a_697_n3946# a_329_n2964# dvdd.t99 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X134 avdd.t395 avdd.t393 avdd.t394 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X135 comparator_0.vpp comparator_0.vpp avdd.t43 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X136 rstring_mux_0.vtrip1.t0 rstring_mux_0.vtrip2.t3 avss.t128 sky130_fd_pr__res_xhigh_po_1p41 l=35
X137 dvss.t695 dvss.t693 osc_ck.t7 dvss.t694 sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X138 comparator_1.vm comparator_1.vm avss.t232 avss.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X139 dvdd.t160 sky130_fd_sc_hd__inv_4_4.Y outb.t12 dvdd.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 avdd.t407 a_429_n1142# a_1636_n1478# avdd.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X141 dvss.t733 a_4653_n2876# a_5860_n3212# dvss.t732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X142 avdd.t89 rstring_mux_0.ena_b rstring_mux_0.vtop.t16 avdd.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X143 avdd.t178 comparator_0.n0 comparator_0.n1 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X144 avdd.t199 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X145 comparator_1.vpp comparator_1.vnn avdd.t147 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X146 dvdd.t103 schmitt_trigger_0.out.t5 schmitt_trigger_0.m.t9 dvdd.t102 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X147 ibias_gen_0.vp0.t11 ibias_gen_0.vp0.t10 avdd.t508 avdd.t507 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X148 outb.t30 sky130_fd_sc_hd__inv_4_4.Y dvss.t415 dvss.t414 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X149 rstring_mux_0.otrip_decoded_avdd[3] a_n4700_n1478# dvss.t555 dvss.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X150 avdd.t392 avdd.t391 avdd.t392 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X151 a_6765_n1142# a_6665_n1230# dvss.t205 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X152 rstring_mux_0.vtop.t15 rstring_mux_0.ena_b avdd.t87 avdd.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X153 ibias_gen_0.ena_b comparator_0.ena avss.t299 avss.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X154 rstring_mux_0.otrip_decoded_avdd[2] a_n4700_n3212# avdd.t111 avdd.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X155 dvdd.t212 otrip_decoded[2].t0 a_n6007_n2964# dvdd.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X156 vin_brout rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.vtrip6.t7 avdd.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X157 avdd.t479 comparator_1.vpp comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X158 avss.t95 avss.t93 avss.t94 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X159 dvss.t89 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t29 dvss.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X160 a_10873_n2760# a_10514_n2760# dvss.t238 dvss.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X161 a_887_n11914# a_509_n19314# avss.t272 sky130_fd_pr__res_xhigh_po_1p41 l=35
X162 comparator_0.vnn comparator_0.vpp avdd.t42 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X163 avdd.t198 comparator_0.vnn comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X164 ibias_gen_0.vp.t4 comparator_0.ena avdd.t558 avdd.t557 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X165 avdd.t485 a_1122_n2256# a_429_n1142# avdd.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X166 osc_ck.t0 rc_osc_0.n.t6 dvss.t146 dvss.t145 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X167 avdd.t85 rstring_mux_0.ena_b rstring_mux_0.vtop.t14 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X168 dvdd.t158 sky130_fd_sc_hd__inv_4_4.Y outb.t11 dvdd.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X169 comparator_0.vt vbg_1v2.t4 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X170 avdd.t93 ibias_gen_0.vp.t8 ibias_gen_0.ibias0 avdd.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X171 dvss.t99 dcomp3v3uv a_10514_n2760# dvss.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X172 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip_decoded_avdd[0] avss.t291 avss.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X173 comparator_1.n1 comparator_1.n0 avss.t361 avss.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X174 ibias_gen_0.vn0.t4 ibias_gen_0.vn0.t3 ibias_gen_0.ve.t4 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X175 ibias_gen_0.vp.t2 ibias_gen_0.isrc_sel_b ibias_gen_0.vp0.t3 avss.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X176 avss.t127 comparator_0.vn comparator_0.vt avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X177 avdd.t390 avdd.t388 avdd.t389 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X178 vin_vunder.t42 avdd.t386 vin_brout avdd.t387 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X179 rstring_mux_0.vtop.t13 rstring_mux_0.ena_b avdd.t83 avdd.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X180 comparator_1.vpp comparator_1.vnn avdd.t146 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X181 ibias_gen_0.vp1.t1 ibias_gen_0.vn1.t10 avss.t145 avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X182 a_n5917_n11914# a_n6295_n19314# avss.t335 sky130_fd_pr__res_xhigh_po_1p41 l=35
X183 avdd.t197 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X184 a_n7751_n2212# a_n8119_n1230# dvss.t670 dvss.t669 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X185 rstring_mux_0.otrip_decoded_avdd[0] a_n6812_n3212# avdd.t216 avdd.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X186 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip_decoded_avdd[4] avss.t218 avss.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X187 dvss.t87 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t28 dvss.t86 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X188 dvss.t627 sky130_fd_sc_hd__inv_4_1.Y vunder.t30 dvss.t626 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X189 dvdd.t235 otrip_decoded[0].t1 a_n8119_n2964# dvdd.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X190 vin_brout rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.vtrip1.t6 avdd.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X191 rc_osc_0.in a_11121_n25357# dvss.t468 sky130_fd_pr__res_xhigh_po_1p41 l=105
X192 dcomp3v3 comparator_1.n1 avdd.t599 avdd.t598 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X193 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvss.t551 dvss.t550 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X194 rstring_mux_0.vtrip_decoded_avdd[1] a_1636_n1478# avdd.t423 avdd.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X195 avdd.t488 a_6765_n1142# a_7972_n1478# avdd.t450 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X196 avdd.t206 a_3234_n2256# a_2541_n1142# avdd.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X197 a_n8195_9395# schmitt_trigger_0.in.t0 avss.t321 sky130_fd_pr__res_xhigh_po_1p41 l=35
X198 rc_osc_0.vr dvdd.t117 rc_osc_0.ena_b dvdd.t118 sky130_fd_pr__pfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.5
X199 vin_brout rstring_mux_0.otrip_decoded_avdd[0] rstring_mux_0.vtrip0.t7 avss.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X200 comparator_0.vnn comparator_0.vpp avdd.t41 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X201 a_n8951_9395# a_n9329_1995# avss.t150 sky130_fd_pr__res_xhigh_po_1p41 l=35
X202 avss.t92 avss.t90 avss.t91 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X203 dcomp.t13 sky130_fd_sc_hd__inv_4_3.Y dvdd.t317 dvdd.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X204 vin_brout avdd.t384 vin_brout avdd.t385 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X205 avdd.t145 comparator_1.vnn comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X206 dvdd.t174 vtrip_decoded[3].t1 a_2441_n1230# dvdd.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X207 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.otrip_decoded_avdd[4] avss.t330 avss.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X208 avdd.t383 avdd.t382 avdd.t383 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X209 vin_vunder.t41 avdd.t380 vin_vunder.t41 avdd.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X210 avdd.t95 ibias_gen_0.vp.t9 itest.t0 avdd.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X211 vin_brout rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.vtrip4.t8 avss.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X212 avdd.t478 comparator_1.vpp comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X213 ibias_gen_0.vstart.t9 vbg_1v2.t5 ibias_gen_0.vn0.t14 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X214 ibias_gen_0.isrc_sel_b avss.t88 ibias_gen_0.ena_b avss.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X215 a_n1683_n1142# a_n1783_n1230# dvss.t118 dvss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X216 comparator_1.vn comparator_0.ena ibias_gen_0.ibias0 avss.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X217 comparator_0.vnn comparator_0.vpp avdd.t40 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X218 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X219 comparator_0.vnn vin_vunder.t51 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X220 a_n20782_n2937# a_n21160_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X221 rstring_mux_0.vtrip_decoded_avdd[3] a_3748_n1478# avdd.t1 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X222 comparator_0.vnn vin_vunder.t52 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X223 dvss.t413 sky130_fd_sc_hd__inv_4_4.Y outb.t29 dvss.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X224 avdd.t415 a_5346_n2256# a_4653_n1142# avdd.t414 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X225 comparator_1.vnn avss.t367 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X226 avdd.t379 avdd.t377 avdd.t378 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X227 comparator_1.vnn avss.t368 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X228 rstring_mux_0.vtop.t12 rstring_mux_0.ena_b avdd.t81 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X229 a_n3795_n1142# a_n3895_n1230# dvss.t263 dvss.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X230 avdd.t144 comparator_1.vnn comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X231 dcomp3v3uv comparator_0.n1 avss.t248 avss.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X232 rstring_mux_0.vtrip5.t6 rstring_mux_0.vtrip_decoded_b_avdd[5] vin_vunder.t20 avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X233 avdd.t447 ibias_gen_0.vp1.t6 ibias_gen_0.vp1.t7 avdd.t446 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X234 vunder.t7 sky130_fd_sc_hd__inv_4_1.Y dvdd.t273 dvdd.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 vin_vunder.t11 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip3.t2 avss.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X236 rc_osc_0.m rc_osc_0.n.t7 dvdd.t59 dvdd.t58 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X237 rstring_mux_0.vtrip3.t8 rstring_mux_0.otrip_decoded_avdd[3] vin_brout avss.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X238 vin_vunder.t29 rstring_mux_0.vtrip_decoded_b_avdd[7] rstring_mux_0.vtrip7.t5 avdd.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X239 avdd.t477 comparator_1.vpp comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X240 dvdd.t233 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvdd.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X241 dvss.t185 a_n6007_n1230# a_n5907_n1142# dvss.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X242 dvss.t532 a_4553_n1230# a_4653_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X243 a_131_n11914# a_n247_n19314# avss.t250 sky130_fd_pr__res_xhigh_po_1p41 l=35
X244 avdd.t376 avdd.t375 avdd.t376 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X245 comparator_1.vn comparator_1.ena_b ibias_gen_0.ibias0 avdd.t524 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X246 avss.t146 ibias_gen_0.vn1.t11 ibias_gen_0.vp1.t2 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X247 avdd.t502 a_7458_n2256# a_6765_n1142# avdd.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X248 rstring_mux_0.vtrip1.t9 rstring_mux_0.vtrip_decoded_avdd[1] vin_vunder.t47 avss.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X249 dvss.t85 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t27 dvss.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X250 avdd.t39 comparator_0.vpp comparator_0.n0 avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X251 rc_osc_0.ena_b osc_ena.t1 dvdd.t132 dvdd.t131 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X252 comparator_0.vt avss.t369 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X253 rstring_mux_0.vtrip0.t6 rstring_mux_0.otrip_decoded_avdd[0] vin_brout avss.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X254 ibias_gen_0.vp1.t3 ibias_gen_0.vn1.t12 avss.t147 avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X255 rstring_mux_0.vtrip_decoded_avdd[6] a_7972_n3212# avdd.t534 avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X256 comparator_0.vnn avss.t370 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X257 avss.t87 avss.t85 avss.t86 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X258 ibias_gen_0.vp.t6 ibias_gen_0.isrc_sel ibias_gen_0.vp0.t7 avdd.t573 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X259 dvss.t728 sky130_fd_sc_hd__inv_4_3.Y dcomp.t30 dvss.t727 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 dvdd.t94 a_10873_n3956# sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X261 dvdd.t156 sky130_fd_sc_hd__inv_4_4.Y outb.t10 dvdd.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X262 vunder.t6 sky130_fd_sc_hd__inv_4_1.Y dvdd.t271 dvdd.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X263 a_n5907_n1142# a_n6007_n1230# dvss.t183 dvss.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X264 comparator_0.n1 comparator_0.n0 avss.t175 avss.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X265 comparator_1.vpp vbg_1v2.t6 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X266 avss.t148 ibias_gen_0.vn1.t13 ibias_gen_0.vp1.t4 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X267 comparator_0.vpp vbg_1v2.t7 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X268 avss.t340 comparator_0.vm comparator_0.vm avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X269 rstring_mux_0.vtrip4.t7 rstring_mux_0.otrip_decoded_avdd[4] vin_brout avss.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X270 dvdd.t237 vtrip_decoded[1].t1 a_329_n1230# dvdd.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X271 a_n10279_n22711# a_11121_n23089# dvss.t698 sky130_fd_pr__res_xhigh_po_1p41 l=105
X272 vin_brout rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.vtrip2.t5 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X273 a_n14999_9395# a_n14621_1995# avss.t263 sky130_fd_pr__res_xhigh_po_1p41 l=35
X274 dcomp3v3uv comparator_0.n1 avdd.t437 avdd.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X275 vin_vunder.t33 rstring_mux_0.vtrip_decoded_b_avdd[3] rstring_mux_0.vtrip3.t5 avdd.t522 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X276 dvdd.t71 vl sky130_fd_sc_hd__inv_4_3.Y dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X277 avdd.t122 a_2541_n1142# a_3748_n1478# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X278 rstring_mux_0.vtrip0.t9 rstring_mux_0.vtrip_decoded_avdd[0] vin_vunder.t38 avss.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X279 rstring_mux_0.vtrip7.t9 rstring_mux_0.otrip_decoded_avdd[7] vin_brout avss.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X280 a_n10463_9395# a_n10085_1995# avss.t195 sky130_fd_pr__res_xhigh_po_1p41 l=35
X281 dvss.t668 a_n8119_n1230# a_n8019_n1142# dvss.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X282 dvss.t204 a_6665_n1230# a_6765_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X283 avdd.t422 a_9570_n2256# a_8877_n1142# avdd.t421 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X284 dvdd.t35 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t13 dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X285 vin_brout avdd.t373 vin_brout avdd.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X286 dvss.t83 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t26 dvss.t82 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X287 dvss.t625 sky130_fd_sc_hd__inv_4_1.Y vunder.t29 dvss.t624 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 comparator_0.vnn comparator_0.vnn avdd.t196 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X289 vin_vunder.t6 avss.t83 vin_vunder.t6 avss.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X290 avdd.t143 comparator_1.vnn comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X291 avdd.t372 avdd.t370 avdd.t372 avdd.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X292 dvss.t639 a_697_n2212# a_1122_n2256# dvss.t638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X293 avdd.t369 avdd.t368 avdd.t369 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X294 a_8877_n1142# a_8777_n1230# dvss.t245 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X295 rc_osc_0.in dvss.t488 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X296 ibias_gen_0.vp.t0 avss.t81 ibias_gen_0.vp.t0 avss.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X297 comparator_1.vn comparator_1.vn avss.t285 avss.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X298 dcomp.t12 sky130_fd_sc_hd__inv_4_3.Y dvdd.t315 dvdd.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 dvss.t13 a_8877_n2876# a_10084_n3212# dvss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X300 a_429_n1142# a_329_n1230# dvss.t544 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X301 rstring_mux_0.otrip_decoded_avdd[6] a_n476_n3212# avdd.t117 avdd.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X302 avdd.t367 avdd.t366 avdd.t367 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X303 a_n11975_9395# a_n12353_1995# avss.t140 sky130_fd_pr__res_xhigh_po_1p41 l=35
X304 avdd.t516 a_4653_n1142# a_5860_n1478# avdd.t515 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X305 dvss.t244 a_8777_n1230# a_8877_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X306 comparator_0.vt vin_vunder.t53 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X307 vin_vunder.t9 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip5.t1 avss.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X308 avdd.t142 comparator_1.vnn comparator_1.vm avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X309 avdd.t219 ibias_gen_0.isrc_sel_b ibias_gen_0.vp0.t4 avdd.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X310 schmitt_trigger_0.m.t4 schmitt_trigger_0.in.t2 dvdd.t83 dvdd.t82 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X311 dvss.t623 sky130_fd_sc_hd__inv_4_1.Y vunder.t28 dvss.t622 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X312 avdd.t365 avdd.t364 avdd.t365 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X313 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.otrip_decoded_avdd[0] avss.t278 avss.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X314 vin_brout avdd.t362 vin_brout avdd.t363 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X315 comparator_1.vnn avss.t371 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X316 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.otrip_decoded_avdd[4] avdd.t580 avdd.t579 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X317 avdd.t361 avdd.t359 avdd.t360 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X318 dvss.t411 sky130_fd_sc_hd__inv_4_4.Y outb.t28 dvss.t410 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X319 a_9203_n11914# a_9581_n19314# avss.t224 sky130_fd_pr__res_xhigh_po_1p41 l=35
X320 dvss.t543 a_329_n1230# a_429_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X321 rc_osc_0.m rc_osc_0.in dvdd.t192 dvdd.t191 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X322 rc_osc_0.m rc_osc_0.in dvss.t487 dvss.t486 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X323 rstring_mux_0.vtrip5.t3 rstring_mux_0.otrip_decoded_avdd[5] vin_brout avss.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X324 avdd.t506 ibias_gen_0.vp0.t8 ibias_gen_0.vp0.t9 avdd.t505 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X325 a_8877_n1142# a_8777_n1230# dvss.t243 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X326 a_n7751_n2212# a_n8119_n1230# dvdd.t289 dvdd.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X327 vin_vunder.t12 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip2.t7 avdd.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X328 avdd.t141 comparator_1.vnn comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X329 rc_osc_0.n.t2 rc_osc_0.m dvdd.t285 dvdd.t284 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X330 a_n6673_n11914# a_n6295_n19314# avss.t123 sky130_fd_pr__res_xhigh_po_1p41 l=35
X331 comparator_0.vt vin_vunder.t54 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X332 avdd.t139 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X333 ibias_gen_0.vn0.t13 vbg_1v2.t8 ibias_gen_0.vstart.t8 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X334 a_5346_n2256# a_4921_n2212# dvss.t680 dvss.t679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X335 avdd.t358 avdd.t356 avdd.t357 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X336 comparator_1.vpp comparator_1.vnn avdd.t138 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X337 avdd.t572 ibias_gen_0.isrc_sel a_n16775_n2223# avdd.t571 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X338 rstring_mux_0.vtrip2.t4 rstring_mux_0.otrip_decoded_avdd[2] vin_brout avss.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X339 dvss.t621 sky130_fd_sc_hd__inv_4_1.Y vunder.t27 dvss.t620 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X340 comparator_1.vm comparator_1.ena_b avss.t270 avss.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X341 dvdd.t231 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvdd.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X342 dcomp3v3 comparator_1.n1 avss.t353 avss.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X343 dvss.t409 sky130_fd_sc_hd__inv_4_4.Y outb.t27 dvss.t408 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X344 avdd.t556 comparator_0.ena ibias_gen_0.vp1.t15 avdd.t555 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X345 avdd.t355 avdd.t354 avdd.t355 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X346 ibias_gen_0.vp1.t17 ibias_gen_0.isrc_sel avdd.t570 avdd.t569 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X347 dcomp.t29 sky130_fd_sc_hd__inv_4_3.Y dvss.t726 dvss.t725 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X348 comparator_0.ena a_10084_n3212# dvss.t356 dvss.t355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X349 rstring_mux_0.vtrip6.t6 rstring_mux_0.otrip_decoded_b_avdd[6] vin_brout avdd.t489 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X350 comparator_1.vpp vbg_1v2.t9 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X351 a_7458_n2256# a_7033_n2212# dvss.t512 dvss.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X352 avdd.t537 a_n1683_n2876# a_n476_n3212# avdd.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X353 rstring_mux_0.vtrip5.t9 rstring_mux_0.vtrip4.t0 avss.t208 sky130_fd_pr__res_xhigh_po_1p41 l=35
X354 comparator_1.vpp vbg_1v2.t10 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X355 vin_vunder.t5 avss.t79 vin_vunder.t5 avss.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X356 sky130_fd_sc_hd__inv_4_3.Y vl dvss.t167 dvss.t166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X357 vunder.t5 sky130_fd_sc_hd__inv_4_1.Y dvdd.t269 dvdd.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X358 avdd.t494 a_n990_n3990# a_n1683_n2876# avdd.t493 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X359 dvdd.t313 sky130_fd_sc_hd__inv_4_3.Y dcomp.t11 dvdd.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X360 brout_filt.t12 sky130_fd_sc_hd__inv_4_0.Y dvdd.t33 dvdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X361 a_n1683_n2876# a_n1783_n2964# dvss.t49 dvss.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X362 dvss.t493 vtrip_decoded[2].t0 a_2441_n2964# dvss.t492 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X363 comparator_0.vn comparator_0.ena_b comparator_0.ibias avdd.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X364 rc_osc_0.in dvss.t485 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X365 a_n9697_n11914# a_n10075_n19314# avss.t211 sky130_fd_pr__res_xhigh_po_1p41 l=35
X366 avss.t246 comparator_0.n1 dcomp3v3uv avss.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X367 avdd.t353 avdd.t352 avdd.t353 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X368 vin_vunder.t4 avss.t77 vin_vunder.t4 avss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X369 comparator_1.vnn comparator_1.vnn avdd.t137 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X370 dvss.t407 sky130_fd_sc_hd__inv_4_4.Y outb.t26 dvss.t406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 comparator_1.vnn comparator_0.ena avdd.t554 avdd.t553 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X372 dcomp3v3 comparator_1.n1 avdd.t597 avdd.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X373 dvss.t81 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t25 dvss.t80 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X374 a_2541_n1142# a_2441_n1230# dvss.t580 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X375 a_n990_n2256# a_n1415_n2212# dvss.t25 dvss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X376 dvdd.t116 dvdd.t114 dvdd.t116 dvdd.t115 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.18
X377 a_n13477_n11914# a_n13099_n19314# avss.t252 sky130_fd_pr__res_xhigh_po_1p41 l=35
X378 dcomp.t28 sky130_fd_sc_hd__inv_4_3.Y dvss.t724 dvss.t723 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X379 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t6 dvdd.t105 dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X380 a_n3795_n1142# a_n3895_n1230# dvss.t261 dvss.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X381 dvss.t731 a_n1683_n1142# a_n476_n1478# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X382 avdd.t457 a_n5214_n2256# a_n5907_n1142# avdd.t456 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X383 rstring_mux_0.vtrip1.t5 rstring_mux_0.otrip_decoded_b_avdd[1] vin_brout avdd.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X384 vin_vunder.t3 avss.t75 vin_vunder.t3 avss.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X385 comparator_0.vn comparator_0.ena_b avss.t171 avss.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X386 ibias_gen_0.vp.t3 avdd.t350 ibias_gen_0.vp.t3 avdd.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X387 a_n10279_n24223# a_11121_n23845# dvss.t382 sky130_fd_pr__res_xhigh_po_1p41 l=105
X388 vunder.t4 sky130_fd_sc_hd__inv_4_1.Y dvdd.t267 dvdd.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X389 dvss.t230 a_n8019_n1142# a_n6812_n1478# dvss.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X390 dvss.t579 a_2441_n1230# a_2541_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X391 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.otrip_decoded_avdd[5] avss.t154 avss.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X392 dcomp3v3uv comparator_0.n1 avss.t244 avss.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X393 avdd.t349 avdd.t348 avdd.t349 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X394 brout_filt.t11 sky130_fd_sc_hd__inv_4_0.Y dvdd.t31 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X395 a_n3795_n2876# a_n3895_n2964# dvss.t37 dvss.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X396 a_2541_n2876# a_2441_n2964# dvss.t574 dvss.t573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X397 comparator_0.vt vin_vunder.t55 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X398 a_n26074_n2937# a_n26452_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X399 a_n23050_n2937# a_n23428_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X400 dvss.t380 a_10515_n2156# a_10874_n2222# dvss.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X401 a_n5161_n11914# a_n4783_n19314# avss.t213 sky130_fd_pr__res_xhigh_po_1p41 l=35
X402 a_n5907_n1142# a_n6007_n1230# dvss.t181 dvss.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X403 rstring_mux_0.vtrip_decoded_avdd[3] a_3748_n1478# dvss.t1 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X404 comparator_0.vnn comparator_0.ena avdd.t552 avdd.t551 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X405 a_n5907_n1142# a_n6007_n1230# dvss.t179 dvss.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X406 a_4653_n1142# a_4553_n1230# dvss.t531 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X407 avdd.t15 a_n7326_n2256# a_n8019_n1142# avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X408 a_n5161_n11914# a_n5539_n19314# avss.t105 sky130_fd_pr__res_xhigh_po_1p41 l=35
X409 avdd.t476 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X410 comparator_1.vnn comparator_1.vnn avdd.t136 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X411 a_n25318_n2937# a_n25696_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X412 ibias_gen_0.vn1.t4 ibias_gen_0.vn1.t3 avss.t144 avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X413 dvss.t253 a_10515_n1026# a_10515_n2156# dvss.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X414 a_n1415_n2212# a_n1783_n1230# dvss.t116 dvss.t115 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X415 dvss.t666 a_n8119_n1230# a_n8019_n1142# dvss.t665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X416 a_4653_n2876# a_4553_n2964# dvss.t290 dvss.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X417 dvss.t269 a_10873_n3956# sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss.t268 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X418 rc_osc_0.in dvss.t484 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X419 avss.t351 comparator_1.n1 dcomp3v3 avss.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X420 a_10873_n3956# a_10514_n3890# dvss.t278 dvss.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X421 a_n8019_n1142# a_n8119_n1230# dvss.t664 dvss.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X422 a_6765_n1142# a_6665_n1230# dvss.t203 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X423 dvss.t491 isrc_sel.t0 a_8777_n1230# dvss.t490 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X424 rstring_mux_0.vtrip2.t1 rstring_mux_0.otrip_decoded_b_avdd[2] vin_brout avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X425 avdd.t347 avdd.t346 avdd.t347 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X426 a_n14999_9395# vl avss.t311 sky130_fd_pr__res_xhigh_po_1p41 l=35
X427 dvss.t619 sky130_fd_sc_hd__inv_4_1.Y vunder.t26 dvss.t618 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X428 a_n8019_n1142# a_n8119_n1230# dvss.t662 dvss.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X429 dvss.t525 vtrip_decoded[0].t0 a_329_n2964# dvss.t524 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X430 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip_decoded_avdd[6] avdd.t531 avdd.t530 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X431 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.otrip_decoded_avdd[7] avss.t364 avss.t363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X432 dvss.t405 sky130_fd_sc_hd__inv_4_4.Y outb.t25 dvss.t404 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 avdd.t38 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X434 a_n3527_n2212# a_n3895_n1230# dvss.t259 dvss.t258 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X435 rstring_mux_0.otrip_decoded_avdd[4] a_n2588_n3212# avdd.t495 avdd.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X436 comparator_1.vnn avss.t372 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X437 a_429_n1142# a_329_n1230# dvss.t542 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X438 a_10873_n2760# a_10514_n2760# dvss.t237 dvss.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X439 dcomp.t27 sky130_fd_sc_hd__inv_4_3.Y dvss.t722 dvss.t721 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X440 vin_vunder.t2 avss.t73 vin_vunder.t2 avss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X441 rstring_mux_0.vtrip2.t6 rstring_mux_0.vtrip_decoded_b_avdd[2] vin_vunder.t13 avdd.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X442 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X443 a_3911_n11914# a_4289_n19314# avss.t109 sky130_fd_pr__res_xhigh_po_1p41 l=35
X444 a_n10463_9395# a_n10841_1995# avss.t287 sky130_fd_pr__res_xhigh_po_1p41 l=35
X445 ibias_gen_0.vp1.t5 ibias_gen_0.vn1.t14 avss.t149 avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X446 a_n8941_n11914# a_n8563_n19314# avss.t256 sky130_fd_pr__res_xhigh_po_1p41 l=35
X447 a_n11965_n11914# a_n11587_n19314# avss.t314 sky130_fd_pr__res_xhigh_po_1p41 l=35
X448 a_6765_n2876# a_6665_n2964# dvss.t593 dvss.t592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X449 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip_decoded_avdd[6] avss.t276 avss.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X450 comparator_0.vt vbg_1v2.t11 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X451 comparator_0.ena_b comparator_0.ena avdd.t550 avdd.t549 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X452 ibias_gen_0.vp0.t5 avdd.t343 avdd.t345 avdd.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X453 avss.t72 avss.t70 avss.t71 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X454 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X455 vunder.t3 sky130_fd_sc_hd__inv_4_1.Y dvdd.t265 dvdd.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 dvss.t465 a_2809_n2212# a_3234_n2256# dvss.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X457 avdd.t342 avdd.t340 avdd.t341 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X458 comparator_1.vnn comparator_1.vnn avdd.t135 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X459 sky130_fd_sc_hd__inv_4_3.Y vl dvss.t165 dvss.t164 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X460 dvss.t541 a_329_n1230# a_429_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X461 dvdd.t206 a_10874_n2222# vl dvdd.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X462 avdd.t475 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X463 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X464 avss.t69 avss.t68 ibias_gen_0.vr.t0 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X465 dvdd.t311 sky130_fd_sc_hd__inv_4_3.Y dcomp.t10 dvdd.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X466 brout_filt.t10 sky130_fd_sc_hd__inv_4_0.Y dvdd.t29 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X467 avss.t242 comparator_0.n1 dcomp3v3uv avss.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X468 dvdd.t154 sky130_fd_sc_hd__inv_4_4.Y outb.t9 dvdd.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X469 avdd.t53 a_8877_n1142# a_10084_n1478# avdd.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X470 avdd.t195 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X471 dvss.t403 sky130_fd_sc_hd__inv_4_4.Y outb.t24 dvss.t402 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X472 a_n5639_n2212# a_n6007_n1230# dvss.t177 dvss.t176 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X473 comparator_0.vpp comparator_0.vpp avdd.t37 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X474 vin_vunder.t39 avdd.t338 vin_vunder.t39 avdd.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X475 a_n9707_9395# a_n9329_1995# avss.t259 sky130_fd_pr__res_xhigh_po_1p41 l=35
X476 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.otrip_decoded_avdd[2] avdd.t107 avdd.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X477 comparator_0.vt vbg_1v2.t12 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X478 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X479 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t7 dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X480 avdd.t36 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X481 dvdd.t41 schmitt_trigger_0.m.t14 schmitt_trigger_0.out.t2 dvdd.t40 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X482 rstring_mux_0.vtop.t11 rstring_mux_0.ena_b avdd.t79 avdd.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X483 vunder.t15 sky130_fd_sc_hd__inv_4_1.Y dvdd.t263 dvdd.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X484 a_n7751_n3946# a_n8119_n2964# dvss.t217 dvss.t216 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X485 a_9570_n2256# a_9145_n2212# dvss.t427 dvss.t426 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X486 dvdd.t309 sky130_fd_sc_hd__inv_4_3.Y dcomp.t9 dvdd.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X487 dvss.t378 a_10515_n2156# a_10874_n2222# dvss.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X488 a_n14989_n11914# a_n15367_n19314# avss.t151 sky130_fd_pr__res_xhigh_po_1p41 l=35
X489 comparator_1.vnn comparator_1.vnn avdd.t134 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X490 comparator_1.n0 comparator_1.ena_b avss.t268 avss.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X491 avdd.t337 avdd.t335 avdd.t337 avdd.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X492 avdd.t443 a_n3795_n2876# a_n2588_n3212# avdd.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X493 a_7458_n2256# a_7033_n2212# dvss.t510 dvss.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X494 a_10514_n3890# a_10514_n2760# avdd.t162 avdd.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X495 a_7691_n11914# a_8069_n19314# avss.t255 sky130_fd_pr__res_xhigh_po_1p41 l=35
X496 dcomp3v3 comparator_1.n1 avss.t349 avss.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X497 a_n10279_n24979# a_11121_n25357# dvss.t168 sky130_fd_pr__res_xhigh_po_1p41 l=105
X498 a_n15745_n11914# a_n15367_n19314# avss.t304 sky130_fd_pr__res_xhigh_po_1p41 l=35
X499 dvss.t114 a_n1783_n1230# a_n1683_n1142# dvss.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X500 dvss.t545 a_4653_n1142# a_5860_n1478# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X501 avdd.t411 a_n3102_n3990# a_n3795_n2876# avdd.t410 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X502 rstring_mux_0.vtrip7.t4 rstring_mux_0.vtrip_decoded_b_avdd[7] vin_vunder.t28 avdd.t491 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X503 avdd.t585 a_n1683_n1142# a_n990_n2256# avdd.t584 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X504 avdd.t334 avdd.t332 avdd.t333 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X505 a_n1683_n2876# a_n1783_n2964# dvss.t47 dvss.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X506 ibias_gen_0.ena_b comparator_0.ena avdd.t548 avdd.t547 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X507 a_n3102_n2256# a_n3527_n2212# dvss.t195 dvss.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X508 avdd.t194 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X509 avdd.t331 avdd.t330 avdd.t331 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X510 comparator_1.vm comparator_1.vnn avdd.t132 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X511 avss.t67 avss.t66 avss.t67 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X512 dvdd.t307 sky130_fd_sc_hd__inv_4_3.Y dcomp.t8 dvdd.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X513 a_2541_n1142# a_2441_n1230# dvss.t578 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X514 ibias_gen_0.isrc_sel a_10084_n1478# avdd.t566 avdd.t565 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X515 dvss.t514 vtrip_decoded[5].t0 a_4553_n1230# dvss.t513 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X516 comparator_0.vpp comparator_0.vpp avdd.t35 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X517 a_2399_n11914# a_2777_n19314# avss.t249 sky130_fd_pr__res_xhigh_po_1p41 l=35
X518 a_10515_n1026# dcomp3v3 avdd.t169 avdd.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X519 avdd.t498 a_n5907_n2876# a_n4700_n3212# avdd.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X520 comparator_0.vt vin_vunder.t56 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X521 ibias_gen_0.vn0.t12 vbg_1v2.t13 ibias_gen_0.vstart.t7 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X522 schmitt_trigger_0.out.t1 schmitt_trigger_0.m.t15 dvdd.t43 dvdd.t42 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X523 a_9570_n2256# a_9145_n2212# dvss.t425 dvss.t424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X524 a_3155_n11914# a_2777_n19314# avss.t214 sky130_fd_pr__res_xhigh_po_1p41 l=35
X525 a_n10453_n11914# a_n10831_n19314# avss.t210 sky130_fd_pr__res_xhigh_po_1p41 l=35
X526 rstring_mux_0.vtrip_decoded_avdd[5] a_5860_n1478# dvss.t558 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X527 dvss.t193 a_n3527_n2212# a_n3102_n2256# dvss.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X528 dvss.t23 a_n1415_n2212# a_n990_n2256# dvss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X529 a_4921_n2212# a_4553_n1230# dvss.t530 dvss.t529 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X530 comparator_1.vnn avss.t373 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X531 dvss.t257 a_n3895_n1230# a_n3795_n1142# dvss.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X532 rstring_mux_0.vtop.t10 rstring_mux_0.ena_b avdd.t77 avdd.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X533 a_n3795_n2876# a_n3895_n2964# dvss.t35 dvss.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X534 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd.t51 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X535 a_n5214_n2256# a_n5639_n2212# dvss.t478 dvss.t477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X536 rstring_mux_0.vtrip_decoded_avdd[4] a_5860_n3212# avdd.t529 avdd.t528 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X537 comparator_0.vt avss.t374 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X538 dvss.t433 vtrip_decoded[7].t0 a_6665_n1230# dvss.t432 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X539 a_131_n11914# a_509_n19314# avss.t129 sky130_fd_pr__res_xhigh_po_1p41 l=35
X540 rc_osc_0.in dvss.t483 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X541 comparator_0.vt vbg_1v2.t14 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X542 avdd.t474 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X543 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X544 a_4653_n1142# a_4553_n1230# dvss.t528 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X545 a_n990_n2256# a_n1415_n2212# dvss.t21 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X546 a_n1415_n2212# a_n1783_n1230# dvdd.t55 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X547 dvss.t134 a_n6007_n2964# a_n5907_n2876# dvss.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X548 dvss.t288 a_4553_n2964# a_4653_n2876# dvss.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X549 outb.t8 sky130_fd_sc_hd__inv_4_4.Y dvdd.t152 dvdd.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 dcomp.t26 sky130_fd_sc_hd__inv_4_3.Y dvss.t720 dvss.t719 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X551 avdd.t418 a_n8019_n2876# a_n6812_n3212# avdd.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X552 ibias_gen_0.vp1.t16 ibias_gen_0.isrc_sel ibias_gen_0.vp.t5 avss.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X553 schmitt_trigger_0.m.t7 schmitt_trigger_0.in.t3 dvss.t219 dvss.t218 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X554 avdd.t329 avdd.t327 avdd.t328 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X555 comparator_0.vpp comparator_0.vpp avdd.t34 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X556 comparator_1.vt avss.t375 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X557 ibias_gen_0.vstart.t6 vbg_1v2.t15 ibias_gen_0.vn0.t11 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X558 dvss.t692 dvss.t690 schmitt_trigger_0.m.t13 dvss.t691 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X559 dvss.t202 a_6665_n1230# a_6765_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X560 rstring_mux_0.vtrip_decoded_avdd[7] a_7972_n1478# dvss.t455 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X561 dvss.t476 a_n5639_n2212# a_n5214_n2256# dvss.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X562 dvss.t482 rc_osc_0.in rc_osc_0.m dvss.t481 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X563 rstring_mux_0.vtop.t9 rstring_mux_0.ena_b avdd.t75 avdd.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X564 avdd.t473 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X565 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X566 dvss.t401 sky130_fd_sc_hd__inv_4_4.Y outb.t23 dvss.t400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X567 dvdd.t190 rc_osc_0.in rc_osc_0.m dvdd.t189 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X568 rc_osc_0.in dvss.t480 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X569 comparator_0.vt avss.t376 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X570 comparator_1.vt avss.t377 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X571 comparator_0.vnn avss.t378 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X572 avss.t339 comparator_0.vm comparator_0.n0 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X573 avdd.t193 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X574 avdd.t326 avdd.t325 avdd.t326 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X575 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X576 sky130_fd_sc_hd__inv_4_4.Y outb_unbuf.t1 dvdd.t176 dvdd.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X577 a_n5907_n2876# a_n6007_n2964# dvss.t132 dvss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X578 dvdd.t198 vtrip_decoded[2].t1 a_2441_n2964# dvdd.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X579 comparator_0.vnn vin_vunder.t57 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X580 ibias_gen_0.isrc_sel_b avdd.t323 ibias_gen_0.ena_b avdd.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X581 brout_filt.t9 sky130_fd_sc_hd__inv_4_0.Y dvdd.t27 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X582 dvdd.t196 isrc_sel.t1 a_8777_n1230# dvdd.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X583 dvdd.t283 rc_osc_0.m rc_osc_0.n.t1 dvdd.t282 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X584 comparator_0.vn comparator_0.vn avss.t126 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X585 a_n7326_n2256# a_n7751_n2212# dvss.t144 dvss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X586 a_6179_n11914# a_6557_n19314# avss.t191 sky130_fd_pr__res_xhigh_po_1p41 l=35
X587 a_n14233_n11914# a_n13855_n19314# avss.t158 sky130_fd_pr__res_xhigh_po_1p41 l=35
X588 comparator_0.vpp vbg_1v2.t16 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X589 avdd.t113 a_429_n2876# a_1636_n3212# avdd.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X590 dvss.t276 a_10514_n3890# a_10873_n3956# dvss.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X591 vin_vunder.t26 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip0.t4 avdd.t420 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X592 a_n23050_n2937# a_n22672_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X593 a_6765_n1142# a_6665_n1230# dvss.t201 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X594 a_n3527_n2212# a_n3895_n1230# dvdd.t91 dvdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X595 comparator_1.vnn comparator_1.vpp avdd.t472 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X596 dvss.t79 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t24 dvss.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X597 dvss.t215 a_n8119_n2964# a_n8019_n2876# dvss.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X598 dvss.t591 a_6665_n2964# a_6765_n2876# dvss.t590 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X599 a_n14233_n11914# a_n14611_n19314# avss.t326 sky130_fd_pr__res_xhigh_po_1p41 l=35
X600 a_n13487_9395# a_n13865_1995# avss.t223 sky130_fd_pr__res_xhigh_po_1p41 l=35
X601 outb.t7 sky130_fd_sc_hd__inv_4_4.Y dvdd.t150 dvdd.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X602 avdd.t322 avdd.t320 avdd.t321 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X603 dvdd.t305 sky130_fd_sc_hd__inv_4_3.Y dcomp.t7 dvdd.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X604 a_1122_n2256# a_697_n2212# dvss.t637 dvss.t636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X605 a_n22294_n2937# a_n21916_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X606 schmitt_trigger_0.m.t3 schmitt_trigger_0.in.t4 dvdd.t85 dvdd.t84 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X607 dvss.t242 a_8777_n1230# a_8877_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X608 dvss.t142 a_n7751_n2212# a_n7326_n2256# dvss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X609 dvss.t446 a_697_n3946# a_1122_n3990# dvss.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X610 rstring_mux_0.vtrip4.t2 rstring_mux_0.otrip_decoded_b_avdd[4] vin_brout avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X611 a_8877_n2876# a_8777_n2964# dvss.t344 dvss.t343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X612 vin_vunder.t32 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip4.t6 avdd.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X613 vunder.t14 sky130_fd_sc_hd__inv_4_1.Y dvdd.t261 dvdd.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X614 avdd.t51 a_8877_n1142# a_9570_n2256# avdd.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X615 dcomp.t25 sky130_fd_sc_hd__inv_4_3.Y dvss.t718 dvss.t717 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X616 avdd.t319 avdd.t317 avdd.t318 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X617 a_1643_n11914# a_1265_n19314# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X618 vin_brout avss.t64 vin_brout avss.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=23.2 ps=169.28 w=5 l=0.6
X619 vunder.t25 sky130_fd_sc_hd__inv_4_1.Y dvss.t617 dvss.t616 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X620 avdd.t5 a_1122_n3990# a_429_n2876# avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X621 comparator_0.n1 comparator_0.n0 avdd.t176 avdd.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X622 avdd.t192 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X623 dvss.t221 schmitt_trigger_0.in.t5 schmitt_trigger_0.m.t6 dvss.t220 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X624 a_429_n2876# a_329_n2964# dvss.t302 dvss.t301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X625 dvss.t549 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvss.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X626 a_8877_n1142# a_8777_n1230# dvss.t241 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X627 a_n5639_n2212# a_n6007_n1230# dvdd.t75 dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X628 dvss.t342 a_8777_n2964# a_8877_n2876# dvss.t341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X629 a_1643_n11914# a_2021_n19314# avss.t310 sky130_fd_pr__res_xhigh_po_1p41 l=35
X630 dvdd.t188 rc_osc_0.in rc_osc_0.m dvdd.t187 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X631 avdd.t316 avdd.t314 avdd.t315 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X632 rstring_mux_0.vtop.t8 rstring_mux_0.ena_b avdd.t73 avdd.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X633 comparator_0.vt vin_vunder.t58 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X634 avss.t63 avss.t60 avss.t62 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X635 dvdd.t303 sky130_fd_sc_hd__inv_4_3.Y dcomp.t6 dvdd.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X636 brout_filt.t8 sky130_fd_sc_hd__inv_4_0.Y dvdd.t25 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X637 a_3234_n2256# a_2809_n2212# dvss.t463 dvss.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X638 rstring_mux_0.vtrip_decoded_b_avdd[1] rstring_mux_0.vtrip_decoded_avdd[1] avdd.t578 avdd.t577 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X639 avss.t313 a_9581_n19314# avss.t312 sky130_fd_pr__res_xhigh_po_1p41 l=35
X640 comparator_0.vt vin_vunder.t59 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X641 avdd.t191 comparator_0.vnn comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X642 comparator_0.vnn comparator_0.vnn avdd.t190 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X643 avdd.t605 comparator_1.n0 comparator_1.n1 avdd.t604 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X644 a_n11219_9395# a_n10841_1995# avss.t309 sky130_fd_pr__res_xhigh_po_1p41 l=35
X645 dvss.t300 a_329_n2964# a_429_n2876# dvss.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X646 avdd.t313 avdd.t311 avdd.t312 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X647 a_8877_n2876# a_8777_n2964# dvss.t340 dvss.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X648 avdd.t71 rstring_mux_0.ena_b rstring_mux_0.vtop.t7 avdd.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X649 comparator_1.vt vbg_1v2.t17 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X650 ibias_gen_0.vp0.t6 comparator_0.ena avdd.t546 avdd.t545 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X651 vin_vunder.t40 avdd.t309 vin_vunder.t40 avdd.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X652 vunder.t24 sky130_fd_sc_hd__inv_4_1.Y dvss.t615 dvss.t614 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X653 rstring_mux_0.vtrip_decoded_avdd[0] a_1636_n3212# avdd.t538 avdd.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X654 avdd.t11 a_6765_n2876# a_7972_n3212# avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X655 avdd.t568 a_3234_n3990# a_2541_n2876# avdd.t567 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X656 rstring_mux_0.vtrip_decoded_b_avdd[5] rstring_mux_0.vtrip_decoded_avdd[5] avdd.t47 avdd.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X657 rstring_mux_0.vtrip_decoded_b_avdd[1] rstring_mux_0.vtrip_decoded_avdd[1] avss.t324 avss.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X658 comparator_1.vnn comparator_1.vpp avdd.t471 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X659 avss.t359 comparator_1.n0 comparator_1.n1 avss.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X660 comparator_1.vt vbg_1v2.t18 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X661 a_5346_n3990# a_4921_n3946# dvss.t649 dvss.t648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X662 ibias_gen_0.vn0.t5 ibias_gen_0.ena_b avss.t166 avss.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X663 dvss.t494 a_6765_n1142# a_7972_n1478# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X664 dvdd.t245 vtrip_decoded[0].t1 a_329_n2964# dvdd.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X665 comparator_0.vt avss.t379 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X666 avss.t240 comparator_0.n1 dcomp3v3uv avss.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X667 a_10515_n2156# a_10515_n1026# avdd.t166 avdd.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X668 rstring_mux_0.vtop.t6 rstring_mux_0.ena_b avdd.t69 avdd.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X669 avdd.t435 comparator_0.n1 dcomp3v3uv avdd.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X670 vin_brout rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.vtrip1.t4 avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X671 a_n10279_n22711# a_11121_n22333# dvss.t169 sky130_fd_pr__res_xhigh_po_1p41 l=105
X672 dcomp3v3 comparator_1.n1 avdd.t595 avdd.t594 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X673 a_n9707_9395# a_n10085_1995# avss.t264 sky130_fd_pr__res_xhigh_po_1p41 l=35
X674 outb.t6 sky130_fd_sc_hd__inv_4_4.Y dvdd.t148 dvdd.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X675 avdd.t520 a_n5907_n1142# a_n5214_n2256# avdd.t519 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X676 dvss.t112 a_n1783_n1230# a_n1683_n1142# dvss.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X677 a_5423_n11914# a_5045_n19314# avss.t194 sky130_fd_pr__res_xhigh_po_1p41 l=35
X678 avdd.t308 avdd.t307 avdd.t308 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X679 avdd.t306 avdd.t304 avdd.t305 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X680 comparator_1.vt avss.t380 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X681 a_n12721_n11914# a_n13099_n19314# avss.t186 sky130_fd_pr__res_xhigh_po_1p41 l=35
X682 comparator_0.vm comparator_0.vnn avdd.t189 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X683 dvss.t163 vl sky130_fd_sc_hd__inv_4_3.Y dvss.t162 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X684 dvdd.t208 vtrip_decoded[5].t1 a_4553_n1230# dvdd.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X685 rstring_mux_0.vtrip_decoded_avdd[2] a_3748_n3212# avdd.t223 avdd.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X686 rstring_mux_0.vtrip3.t9 rstring_mux_0.vtrip4.t9 avss.t336 sky130_fd_pr__res_xhigh_po_1p41 l=35
X687 avdd.t225 a_5346_n3990# a_4653_n2876# avdd.t224 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X688 a_7458_n3990# a_7033_n3946# dvss.t350 dvss.t349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X689 schmitt_trigger_0.in.t6 dvss.t222 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X690 vunder.t13 sky130_fd_sc_hd__inv_4_1.Y dvdd.t259 dvdd.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X691 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.otrip_decoded_avdd[3] avss.t333 avss.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X692 vin_brout avdd.t302 vin_brout avdd.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X693 sky130_fd_sc_hd__inv_4_4.Y outb_unbuf.t2 dvdd.t178 dvdd.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X694 rstring_mux_0.vtrip3.t0 rstring_mux_0.vtrip2.t2 avss.t103 sky130_fd_pr__res_xhigh_po_1p41 l=35
X695 avss.t59 avss.t57 avss.t58 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X696 a_n1683_n1142# a_n1783_n1230# dvss.t110 dvss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X697 rc_osc_0.m rc_osc_0.n.t8 dvdd.t61 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X698 vin_brout avss.t55 vin_brout avss.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X699 comparator_1.ena_b comparator_0.ena avss.t296 avss.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X700 avdd.t301 avdd.t300 avdd.t301 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X701 brout_filt.t23 sky130_fd_sc_hd__inv_4_0.Y dvss.t77 dvss.t76 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X702 a_4921_n2212# a_4553_n1230# dvdd.t218 dvdd.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X703 dcomp3v3uv comparator_0.n1 avdd.t433 avdd.t432 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X704 comparator_0.vnn comparator_0.vnn avdd.t188 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X705 avdd.t299 avdd.t297 avdd.t298 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X706 a_9570_n2256# a_9145_n2212# dvss.t423 dvss.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X707 dvss.t274 a_10514_n3890# a_10873_n3956# dvss.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X708 dvdd.t109 schmitt_trigger_0.out.t8 sky130_fd_sc_hd__inv_4_0.Y dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X709 comparator_0.vt vbg_1v2.t19 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X710 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X711 dvss.t577 a_2441_n1230# a_2541_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X712 dvss.t19 a_n1415_n2212# a_n990_n2256# dvss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X713 schmitt_trigger_0.in.t7 dvss.t223 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X714 avdd.t131 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X715 ibias_gen_0.vn1.t0 avss.t53 ibias_gen_0.vp1.t0 avss.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X716 dcomp.t24 sky130_fd_sc_hd__inv_4_3.Y dvss.t716 dvss.t715 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X717 avdd.t160 a_n8019_n1142# a_n7326_n2256# avdd.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X718 dvss.t255 a_n3895_n1230# a_n3795_n1142# dvss.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X719 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t9 dvss.t304 dvss.t303 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X720 dvdd.t257 sky130_fd_sc_hd__inv_4_1.Y vunder.t12 dvdd.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X721 a_2541_n2876# a_2441_n2964# dvss.t572 dvss.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X722 a_n990_n3990# a_n1415_n3946# dvss.t61 dvss.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X723 avdd.t296 avdd.t294 avdd.t295 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X724 vin_vunder.t36 rstring_mux_0.vtrip_decoded_avdd[6] rstring_mux_0.vtrip6.t9 avss.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X725 ibias_gen_0.vn0.t10 vbg_1v2.t20 ibias_gen_0.vstart.t5 avss.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X726 dvdd.t172 vtrip_decoded[7].t1 a_6665_n1230# dvdd.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X727 a_n3795_n2876# a_n3895_n2964# dvss.t33 dvss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X728 dvss.t557 a_n5907_n1142# a_n4700_n1478# dvss.t556 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X729 a_n5214_n2256# a_n5639_n2212# dvss.t474 dvss.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X730 a_n7751_n3946# a_n8119_n2964# dvdd.t79 dvdd.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X731 avdd.t527 a_7458_n3990# a_6765_n2876# avdd.t526 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X732 rc_osc_0.vr dvss.t687 dvss.t689 dvss.t688 sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X733 avdd.t32 comparator_0.vpp comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X734 a_n3102_n2256# a_n3527_n2212# dvss.t191 dvss.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X735 a_n990_n2256# a_n1415_n2212# dvss.t17 dvss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X736 dvss.t502 a_10874_n2222# vl dvss.t501 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X737 avss.t230 comparator_1.vm comparator_1.n0 avss.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X738 dvdd.t87 schmitt_trigger_0.in.t8 schmitt_trigger_0.m.t2 dvdd.t86 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X739 brout_filt.t7 sky130_fd_sc_hd__inv_4_0.Y dvdd.t23 dvdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X740 vin_brout rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.vtrip2.t0 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X741 a_8447_n11914# a_8825_n19314# avss.t220 sky130_fd_pr__res_xhigh_po_1p41 l=35
X742 brout_filt.t22 sky130_fd_sc_hd__inv_4_0.Y dvss.t75 dvss.t74 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X743 rstring_mux_0.vtrip_decoded_avdd[1] a_1636_n1478# dvss.t434 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X744 dvss.t570 a_2441_n2964# a_2541_n2876# dvss.t569 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X745 rstring_mux_0.vtrip0.t3 rstring_mux_0.vtrip_decoded_b_avdd[0] vin_vunder.t25 avdd.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X746 a_10873_n2760# a_10873_n3956# dvdd.t93 dvdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X747 rstring_mux_0.vtrip0.t2 rstring_mux_0.otrip_decoded_b_avdd[0] vin_brout avdd.t413 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X748 dvss.t547 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvss.t546 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 a_9203_n11914# a_8825_n19314# avss.t139 sky130_fd_pr__res_xhigh_po_1p41 l=35
X750 dvss.t175 a_n6007_n1230# a_n5907_n1142# dvss.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X751 a_n5917_n11914# a_n5539_n19314# avss.t251 sky130_fd_pr__res_xhigh_po_1p41 l=35
X752 comparator_0.vnn comparator_0.vnn avdd.t187 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X753 rstring_mux_0.vtrip7.t7 rstring_mux_0.vtrip_decoded_avdd[7] vin_vunder.t45 avss.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X754 a_n5907_n2876# a_n6007_n2964# dvss.t130 dvss.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X755 avdd.t293 avdd.t291 avdd.t292 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X756 a_n5907_n2876# a_n6007_n2964# dvss.t128 dvss.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X757 a_4653_n2876# a_4553_n2964# dvss.t286 dvss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X758 comparator_0.n0 comparator_0.ena_b avss.t169 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X759 avdd.t290 avdd.t289 avdd.t290 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X760 dvdd.t301 sky130_fd_sc_hd__inv_4_3.Y dcomp.t5 dvdd.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X761 avdd.t55 a_2541_n2876# a_3748_n3212# avdd.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X762 avss.t121 rstring_mux_0.ena_b rstring_mux_0.vtop.t0 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X763 avdd.t130 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X764 avss.t260 ibias_gen_0.vn1.t15 ibias_gen_0.vp1.t12 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X765 a_n7326_n2256# a_n7751_n2212# dvss.t140 dvss.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X766 avdd.t103 a_9570_n3990# a_8877_n2876# avdd.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X767 vin_brout rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.vtrip3.t7 avss.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X768 rstring_mux_0.vtrip4.t5 rstring_mux_0.vtrip_decoded_b_avdd[4] vin_vunder.t31 avdd.t503 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X769 comparator_1.vnn comparator_1.vpp avdd.t470 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X770 comparator_1.vt vbg_1v2.t21 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X771 a_n8019_n1142# a_n8119_n1230# dvss.t660 dvss.t659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X772 a_n1415_n3946# a_n1783_n2964# dvss.t45 dvss.t44 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X773 comparator_0.vt comparator_0.vn avss.t125 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X774 ibias_gen_0.vstart.t4 vbg_1v2.t22 ibias_gen_0.vn0.t9 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X775 dvss.t213 a_n8119_n2964# a_n8019_n2876# dvss.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X776 vin_vunder.t1 avss.t51 vin_vunder.t1 avss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X777 vunder.t23 sky130_fd_sc_hd__inv_4_1.Y dvss.t613 dvss.t612 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X778 a_3911_n11914# a_3533_n19314# avss.t341 sky130_fd_pr__res_xhigh_po_1p41 l=35
X779 vin_brout rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.vtrip6.t4 avss.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X780 a_1122_n2256# a_697_n2212# dvss.t635 dvss.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X781 dvss.t272 a_10514_n3890# a_10873_n3956# dvss.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X782 comparator_1.vnn comparator_1.vpp avdd.t469 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X783 avss.t50 avss.t48 avss.t49 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X784 a_10874_n1026# a_10515_n1026# dvss.t251 dvss.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X785 a_n8019_n2876# a_n8119_n2964# dvss.t211 dvss.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X786 a_6765_n2876# a_6665_n2964# dvss.t589 dvss.t588 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X787 dvss.t373 ena.t0 a_8777_n2964# dvss.t372 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X788 comparator_0.ibias ibias_gen_0.vp.t10 avdd.t97 avdd.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X789 dvss.t461 a_2809_n2212# a_3234_n2256# dvss.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X790 a_n8019_n2876# a_n8119_n2964# dvss.t209 dvss.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X791 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.otrip_decoded_avdd[0] avdd.t533 avdd.t532 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X792 dvdd.t49 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X sky130_fd_sc_hd__inv_4_1.A dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X793 avdd.t606 a_4653_n2876# a_5860_n3212# avdd.t528 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X794 dvss.t236 a_10514_n2760# a_10873_n2760# dvss.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X795 rstring_mux_0.vtrip5.t8 rstring_mux_0.vtrip6.t5 avss.t192 sky130_fd_pr__res_xhigh_po_1p41 l=35
X796 osc_ck.t3 rc_osc_0.ena_b rc_osc_0.vr dvdd.t95 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X797 dvss.t267 dcomp3v3 a_10515_n1026# dvss.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X798 dvss.t633 a_697_n2212# a_1122_n2256# dvss.t632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X799 a_n3527_n3946# a_n3895_n2964# dvss.t31 dvss.t30 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X800 a_429_n2876# a_329_n2964# dvss.t298 dvss.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X801 vin_brout rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.vtrip7.t8 avss.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X802 dvss.t385 osc_ena.t2 rc_osc_0.ena_b dvss.t384 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X803 a_n14243_9395# a_n13865_1995# avss.t207 sky130_fd_pr__res_xhigh_po_1p41 l=35
X804 vunder.t22 sky130_fd_sc_hd__inv_4_1.Y dvss.t611 dvss.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X805 vin_vunder.t22 rstring_mux_0.vtrip_decoded_avdd[4] rstring_mux_0.vtrip4.t3 avss.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X806 avdd.t468 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X807 outb.t5 sky130_fd_sc_hd__inv_4_4.Y dvdd.t146 dvdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X808 a_3234_n2256# a_2809_n2212# dvss.t459 dvss.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X809 rstring_mux_0.vtrip7.t0 rstring_mux_0.vtrip6.t0 avss.t102 sky130_fd_pr__res_xhigh_po_1p41 l=35
X810 a_n9697_n11914# a_n9319_n19314# avss.t98 sky130_fd_pr__res_xhigh_po_1p41 l=35
X811 avdd.t288 avdd.t287 avdd.t288 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X812 comparator_0.vt vbg_1v2.t23 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X813 schmitt_trigger_0.out.t0 schmitt_trigger_0.m.t16 dvdd.t45 dvdd.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X814 avdd.t453 a_n3795_n1142# a_n3102_n2256# avdd.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X815 dvss.t320 a_2809_n3946# a_3234_n3990# dvss.t319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X816 a_n10279_n23467# a_11121_n23845# dvss.t159 sky130_fd_pr__res_xhigh_po_1p41 l=105
X817 comparator_1.vn comparator_1.ena_b avss.t266 avss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X818 brout_filt.t21 sky130_fd_sc_hd__inv_4_0.Y dvss.t73 dvss.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X819 dvss.t296 a_329_n2964# a_429_n2876# dvss.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X820 comparator_0.vt avss.t381 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X821 comparator_0.vt vbg_1v2.t24 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X822 avdd.t31 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X823 dvss.t399 sky130_fd_sc_hd__inv_4_4.Y outb.t22 dvss.t398 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X824 rstring_mux_0.otrip_decoded_avdd[7] a_n476_n1478# dvss.t270 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X825 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X826 dvss.t678 a_4921_n2212# a_5346_n2256# dvss.t677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X827 vin_vunder.t44 rstring_mux_0.vtrip_decoded_avdd[7] rstring_mux_0.vtrip7.t6 avss.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X828 avdd.t593 comparator_1.n1 dcomp3v3 avdd.t592 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X829 avss.t209 a_n27208_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X830 a_n5639_n3946# a_n6007_n2964# dvss.t126 dvss.t125 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X831 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t10 dvss.t306 dvss.t305 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 dvdd.t255 sky130_fd_sc_hd__inv_4_1.Y vunder.t11 dvdd.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X833 rstring_mux_0.vtrip5.t0 rstring_mux_0.vtrip_decoded_avdd[5] vin_vunder.t8 avss.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X834 comparator_1.vt avss.t382 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X835 ibias_gen_0.ibias0 ibias_gen_0.vp.t11 avdd.t99 avdd.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X836 rstring_mux_0.vtrip5.t5 rstring_mux_0.otrip_decoded_b_avdd[5] vin_brout avdd.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X837 a_5346_n2256# a_4921_n2212# dvss.t676 dvss.t675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X838 rstring_mux_0.vtrip_decoded_b_avdd[3] rstring_mux_0.vtrip_decoded_avdd[3] avdd.t105 avdd.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X839 a_n4405_n11914# a_n4783_n19314# avss.t258 sky130_fd_pr__res_xhigh_po_1p41 l=35
X840 avss.t238 comparator_0.n1 dcomp3v3uv avss.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X841 comparator_0.vpp comparator_0.ena avdd.t544 avdd.t543 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X842 vin_brout rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.vtrip5.t2 avss.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X843 avdd.t286 avdd.t284 avdd.t285 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X844 a_9570_n3990# a_9145_n3946# dvss.t156 dvss.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X845 avdd.t467 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X846 avss.t47 avss.t46 avss.t47 avss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X847 avdd.t405 a_429_n1142# a_1122_n2256# avdd.t404 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X848 avdd.t283 avdd.t282 avdd.t283 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X849 comparator_1.vnn avss.t383 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X850 dvss.t508 a_7033_n2212# a_7458_n2256# dvss.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X851 avdd.t431 comparator_0.n1 dcomp3v3uv avdd.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X852 a_n15479_n3901# ibias_gen_0.isrc_sel ibias_gen_0.vn1.t9 avss.t319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X853 dcomp.t23 sky130_fd_sc_hd__inv_4_3.Y dvss.t714 dvss.t713 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X854 dvss.t224 a_2541_n1142# a_3748_n1478# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X855 outb.t4 sky130_fd_sc_hd__inv_4_4.Y dvdd.t144 dvdd.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X856 rstring_mux_0.otrip_decoded_avdd[2] a_n4700_n3212# dvss.t171 dvss.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X857 a_7458_n3990# a_7033_n3946# dvss.t348 dvss.t347 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X858 rstring_mux_0.vtrip_decoded_b_avdd[3] rstring_mux_0.vtrip_decoded_avdd[3] avss.t133 avss.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X859 comparator_0.n0 comparator_0.vpp avdd.t30 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X860 avdd.t591 comparator_1.n1 dcomp3v3 avdd.t590 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X861 schmitt_trigger_0.m.t10 schmitt_trigger_0.out.t11 dvdd.t111 dvdd.t110 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X862 dvdd.t63 rc_osc_0.n.t9 osc_ck.t1 dvdd.t62 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X863 rc_osc_0.m rc_osc_0.n.t10 dvss.t148 dvss.t147 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X864 dvss.t43 a_n1783_n2964# a_n1683_n2876# dvss.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X865 avss.t45 avss.t44 avss.t45 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X866 ibias_gen_0.vp0.t1 ibias_gen_0.vn0.t20 ibias_gen_0.vr.t2 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X867 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss.t106 dvss.t105 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X868 a_2809_n2212# a_2441_n1230# dvss.t576 dvss.t575 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X869 avdd.t29 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X870 brout_filt.t6 sky130_fd_sc_hd__inv_4_0.Y dvdd.t21 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X871 dvss.t189 a_n3527_n2212# a_n3102_n2256# dvss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X872 avdd.t483 a_n5214_n3990# a_n5907_n2876# avdd.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X873 vunder.t21 sky130_fd_sc_hd__inv_4_1.Y dvss.t609 dvss.t608 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X874 a_n3102_n3990# a_n3527_n3946# dvss.t330 dvss.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X875 a_2541_n2876# a_2441_n2964# dvss.t568 dvss.t567 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X876 dvss.t431 vtrip_decoded[4].t0 a_4553_n2964# dvss.t430 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X877 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.otrip_decoded_avdd[5] avdd.t119 avdd.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X878 avdd.t121 a_2541_n1142# a_3234_n2256# avdd.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X879 dvss.t421 a_9145_n2212# a_9570_n2256# dvss.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X880 rstring_mux_0.vtrip7.t3 rstring_mux_0.otrip_decoded_b_avdd[7] vin_brout avdd.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X881 dcomp3v3 comparator_1.n1 avss.t347 avss.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X882 a_n8185_n11914# a_n7807_n19314# avss.t271 sky130_fd_pr__res_xhigh_po_1p41 l=35
X883 vin_vunder.t18 rstring_mux_0.vtrip_decoded_avdd[2] rstring_mux_0.vtrip2.t8 avss.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X884 a_n3102_n2256# a_n3527_n2212# dvss.t187 dvss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X885 rstring_mux_0.otrip_decoded_avdd[0] a_n6812_n3212# dvss.t332 dvss.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X886 a_9570_n3990# a_9145_n3946# dvss.t154 dvss.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X887 dvss.t328 a_n3527_n3946# a_n3102_n3990# dvss.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X888 dvss.t59 a_n1415_n3946# a_n990_n3990# dvss.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X889 a_4921_n3946# a_4553_n2964# dvss.t284 dvss.t283 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X890 comparator_1.vpp comparator_1.vpp avdd.t466 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X891 dvss.t29 a_n3895_n2964# a_n3795_n2876# dvss.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X892 dvss.t234 a_10514_n2760# a_10873_n2760# dvss.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X893 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip_decoded_avdd[2] avdd.t158 avdd.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X894 a_n11209_n11914# a_n11587_n19314# avss.t212 sky130_fd_pr__res_xhigh_po_1p41 l=35
X895 comparator_0.vpp comparator_0.vnn avdd.t186 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X896 vin_vunder.t27 avdd.t280 vin_vunder.t27 avdd.t281 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X897 avdd.t279 avdd.t277 avdd.t278 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X898 schmitt_trigger_0.m.t11 schmitt_trigger_0.out.t12 dvss.t308 dvss.t307 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X899 comparator_0.ena_b comparator_0.ena avss.t294 avss.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X900 a_7033_n2212# a_6665_n1230# dvss.t199 dvss.t198 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X901 comparator_1.vt vbg_1v2.t25 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X902 dvss.t472 a_n5639_n2212# a_n5214_n2256# dvss.t471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X903 avdd.t17 a_n7326_n3990# a_n8019_n2876# avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X904 dvss.t527 a_4553_n1230# a_4653_n1142# dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X905 a_n5214_n3990# a_n5639_n3946# dvss.t368 dvss.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X906 avss.t284 comparator_1.vn comparator_1.vt avss.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X907 dvss.t371 otrip_decoded[7].t0 a_n1783_n1230# dvss.t370 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X908 dvss.t522 vtrip_decoded[6].t0 a_6665_n2964# dvss.t521 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X909 comparator_0.vt avss.t384 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X910 vunder.t20 sky130_fd_sc_hd__inv_4_1.Y dvss.t607 dvss.t606 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X911 avdd.t514 a_4653_n1142# a_5346_n2256# avdd.t513 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X912 a_4653_n2876# a_4553_n2964# dvss.t282 dvss.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X913 a_n990_n3990# a_n1415_n3946# dvss.t57 dvss.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X914 comparator_0.vnn avss.t385 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X915 vin_brout rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.vtrip4.t1 avdd.t402 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X916 outb.t21 sky130_fd_sc_hd__inv_4_4.Y dvss.t397 dvss.t396 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X917 comparator_0.vt avss.t386 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X918 comparator_0.vpp vbg_1v2.t26 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X919 vin_vunder.t17 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip6.t2 avdd.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X920 comparator_1.n0 comparator_1.vm avss.t228 avss.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X921 dvdd.t180 outb_unbuf.t3 sky130_fd_sc_hd__inv_4_4.Y dvdd.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X922 a_n5214_n2256# a_n5639_n2212# dvss.t470 dvss.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X923 dvss.t587 a_6665_n2964# a_6765_n2876# dvss.t586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X924 dvss.t366 a_n5639_n3946# a_n5214_n3990# dvss.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X925 avdd.t28 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X926 sky130_fd_sc_hd__inv_4_4.Y outb_unbuf.t4 dvss.t450 dvss.t449 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X927 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.otrip_decoded_avdd[7] avdd.t610 avdd.t609 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X928 avdd.t276 avdd.t275 avdd.t276 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X929 comparator_1.vt avss.t387 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X930 brout_filt.t20 sky130_fd_sc_hd__inv_4_0.Y dvss.t71 dvss.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X931 a_1122_n2256# a_697_n2212# dvss.t631 dvss.t630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X932 a_9145_n2212# a_8777_n1230# dvss.t240 dvss.t239 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X933 comparator_0.vnn avss.t388 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X934 dvss.t138 a_n7751_n2212# a_n7326_n2256# dvss.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X935 comparator_0.vnn vin_vunder.t60 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X936 comparator_1.vpp comparator_1.vpp avdd.t465 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X937 dvss.t161 vl sky130_fd_sc_hd__inv_4_3.Y dvss.t160 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X938 a_n7326_n3990# a_n7751_n3946# dvss.t9 dvss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X939 comparator_0.vpp comparator_0.vnn avdd.t185 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X940 dvss.t520 otrip_decoded[5].t0 a_n3895_n1230# dvss.t519 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X941 comparator_0.vpp vbg_1v2.t27 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X942 outb.t3 sky130_fd_sc_hd__inv_4_4.Y dvdd.t142 dvdd.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X943 avdd.t487 a_6765_n1142# a_7458_n2256# avdd.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X944 a_6765_n2876# a_6665_n2964# dvss.t585 dvss.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X945 comparator_1.vnn avss.t389 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X946 outb.t20 sky130_fd_sc_hd__inv_4_4.Y dvss.t395 dvss.t394 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X947 a_697_n2212# a_329_n1230# dvss.t540 dvss.t539 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X948 avdd.t464 comparator_1.vpp comparator_1.vnn avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X949 comparator_1.vnn avss.t390 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X950 a_1122_n3990# a_697_n3946# dvss.t444 dvss.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X951 a_n26074_n2937# a_n25696_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X952 avdd.t274 avdd.t273 avdd.t274 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X953 dvdd.t113 schmitt_trigger_0.out.t13 sky130_fd_sc_hd__inv_4_0.Y dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X954 dvss.t338 a_8777_n2964# a_8877_n2876# dvss.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X955 dvss.t7 a_n7751_n3946# a_n7326_n3990# dvss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X956 a_n11219_9395# a_n11597_1995# avss.t106 sky130_fd_pr__res_xhigh_po_1p41 l=35
X957 dcomp.t22 sky130_fd_sc_hd__inv_4_3.Y dvss.t712 dvss.t711 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X958 avss.t345 comparator_1.n1 dcomp3v3 avss.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X959 rstring_mux_0.vtrip_decoded_b_avdd[7] rstring_mux_0.vtrip_decoded_avdd[7] avdd.t564 avdd.t563 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X960 a_n12731_9395# a_n12353_1995# avss.t107 sky130_fd_pr__res_xhigh_po_1p41 l=35
X961 a_429_n1142# a_329_n1230# dvss.t538 dvss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X962 a_3234_n2256# a_2809_n2212# dvss.t457 dvss.t456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X963 a_n25318_n2937# a_n24940_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X964 avdd.t9 a_8877_n2876# a_10084_n3212# avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X965 avdd.t27 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X966 avdd.t272 avdd.t271 avdd.t272 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X967 rstring_mux_0.vtrip_decoded_avdd[6] a_7972_n3212# dvss.t562 dvss.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X968 vin_brout rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.vtrip5.t4 avdd.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X969 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss.t104 dvss.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X970 dvss.t496 otrip_decoded[3].t0 a_n6007_n1230# dvss.t495 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X971 a_8877_n2876# a_8777_n2964# dvss.t336 dvss.t335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X972 osc_ck.t2 rc_osc_0.n.t11 dvdd.t65 dvdd.t64 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X973 avss.t318 ibias_gen_0.isrc_sel ibias_gen_0.vn0.t18 avss.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X974 dvdd.t299 sky130_fd_sc_hd__inv_4_3.Y dcomp.t4 dvdd.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X975 brout_filt.t5 sky130_fd_sc_hd__inv_4_0.Y dvdd.t19 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X976 dvss.t674 a_4921_n2212# a_5346_n2256# dvss.t673 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X977 avss.t316 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b avss.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X978 brout_filt.t19 sky130_fd_sc_hd__inv_4_0.Y dvss.t69 dvss.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X979 a_n1415_n3946# a_n1783_n2964# dvdd.t3 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X980 a_3234_n3990# a_2809_n3946# dvss.t318 dvss.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X981 a_7691_n11914# a_7313_n19314# avss.t253 sky130_fd_pr__res_xhigh_po_1p41 l=35
X982 avdd.t26 comparator_0.vpp comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X983 comparator_1.vpp comparator_1.vpp avdd.t463 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X984 a_n22294_n2937# a_n22672_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X985 a_5346_n2256# a_4921_n2212# dvss.t672 dvss.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X986 comparator_1.vnn comparator_1.vpp avdd.t462 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X987 ibias_gen_0.vp1.t10 ibias_gen_0.isrc_sel_b ibias_gen_0.vp.t1 avdd.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X988 avdd.t67 rstring_mux_0.ena_b rstring_mux_0.vtop.t5 avdd.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X989 dvss.t500 otrip_decoded[1].t0 a_n8119_n1230# dvss.t499 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X990 comparator_1.vt vbg_1v2.t28 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X991 dvdd.t168 ena.t1 a_8777_n2964# dvdd.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X992 dvss.t686 dvss.t684 rc_osc_0.m dvss.t685 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X993 a_n24562_n2937# a_n24940_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X994 a_n21538_n2937# a_n21916_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X995 dvss.t506 a_7033_n2212# a_7458_n2256# dvss.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X996 dvdd.t221 rc_osc_0.n.t12 rc_osc_0.m dvdd.t220 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X997 comparator_1.vpp vbg_1v2.t29 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X998 a_n3527_n3946# a_n3895_n2964# dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X999 comparator_0.vnn avss.t391 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1000 ibias_gen_0.vstart.t3 vbg_1v2.t30 ibias_gen_0.vn0.t8 avss.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1001 avss.t142 ibias_gen_0.vn1.t1 ibias_gen_0.vn1.t2 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1002 rstring_mux_0.otrip_decoded_avdd[6] a_n476_n3212# dvss.t197 dvss.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1003 avdd.t536 a_n1683_n2876# a_n990_n3990# avdd.t535 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1004 vin_brout rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.vtrip7.t2 avdd.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1005 comparator_1.vpp vbg_1v2.t31 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1006 outb.t19 sky130_fd_sc_hd__inv_4_4.Y dvss.t393 dvss.t392 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1007 a_n10279_n24979# a_11121_n24601# dvss.t489 sky130_fd_pr__res_xhigh_po_1p41 l=105
X1008 avdd.t129 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1009 avss.t41 avss.t39 avss.t41 avss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1010 a_n23806_n2937# a_n24184_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1011 avss.t164 ibias_gen_0.ena_b ibias_gen_0.vn1.t5 avss.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1012 a_2809_n2212# a_2441_n1230# dvdd.t241 dvdd.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1013 dvss.t41 a_n1783_n2964# a_n1683_n2876# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1014 comparator_0.vpp vbg_1v2.t32 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1015 vunder.t19 sky130_fd_sc_hd__inv_4_1.Y dvss.t605 dvss.t604 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 a_7458_n2256# a_7033_n2212# dvss.t504 dvss.t503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1017 comparator_0.ena a_10084_n3212# avdd.t222 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1018 rc_osc_0.vr a_11121_n22333# dvss.t369 sky130_fd_pr__res_xhigh_po_1p41 l=105
X1019 avdd.t65 rstring_mux_0.ena_b rstring_mux_0.vtop.t4 avdd.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1020 dcomp3v3 comparator_1.n1 avss.t343 avss.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1021 dvdd.t47 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X sky130_fd_sc_hd__inv_4_1.A dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1022 rstring_mux_0.vtrip_decoded_b_avdd[5] rstring_mux_0.vtrip_decoded_avdd[5] avss.t111 avss.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1023 comparator_1.vpp comparator_1.vpp avdd.t461 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1024 sky130_fd_sc_hd__inv_4_4.Y outb_unbuf.t5 dvss.t452 dvss.t451 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1025 vin_brout rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.vtrip0.t1 avdd.t412 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1026 comparator_0.vm comparator_0.vm avss.t338 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1027 avss.t43 avss.t42 ibias_gen_0.ve.t1 avss sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544 d=4547244,10712
X1028 ibias_gen_0.isrc_sel a_10084_n1478# dvss.t658 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1029 comparator_0.vt vin_vunder.t61 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1030 comparator_1.vnn comparator_1.vpp avdd.t460 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1031 avss.t38 avss.t37 avss.t38 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1032 dvss.t710 sky130_fd_sc_hd__inv_4_3.Y dcomp.t21 dvss.t709 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1033 dvdd.t279 schmitt_trigger_0.in.t9 schmitt_trigger_0.m.t1 dvdd.t278 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1034 dvss.t419 a_9145_n2212# a_9570_n2256# dvss.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1035 a_n1683_n2876# a_n1783_n2964# dvss.t39 dvss.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1036 ibias_gen_0.ve.t0 avss.t35 avss.t36 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1037 schmitt_trigger_0.m.t0 schmitt_trigger_0.in.t10 dvdd.t281 dvdd.t280 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1038 rstring_mux_0.otrip_decoded_avdd[3] a_n4700_n1478# avdd.t518 avdd.t517 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1039 a_n5639_n3946# a_n6007_n2964# dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1040 avdd.t429 comparator_0.n1 dcomp3v3uv avdd.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1041 dvss.t516 schmitt_trigger_0.out.t14 sky130_fd_sc_hd__inv_4_0.Y dvss.t515 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1042 a_9570_n3990# a_9145_n3946# dvss.t152 dvss.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1043 dvdd.t253 sky130_fd_sc_hd__inv_4_1.Y vunder.t10 dvdd.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1044 a_7033_n2212# a_6665_n1230# dvdd.t77 dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1045 dvss.t566 a_2441_n2964# a_2541_n2876# dvss.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1046 dvss.t55 a_n1415_n3946# a_n990_n3990# dvss.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1047 a_n8185_n11914# a_n8563_n19314# avss.t254 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1048 dvss.t27 a_n3895_n2964# a_n3795_n2876# dvss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1049 rstring_mux_0.vtrip6.t1 rstring_mux_0.vtrip_decoded_b_avdd[6] vin_vunder.t16 avdd.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1050 ibias_gen_0.vp1.t13 ibias_gen_0.vn1.t16 avss.t261 avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1051 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvdd.t229 dvdd.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1052 dvss.t467 a_n3795_n1142# a_n2588_n1478# dvss.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1053 avss.t262 ibias_gen_0.vn1.t17 ibias_gen_0.vp1.t14 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1054 dvdd.t17 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t4 dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1055 dvdd.t130 otrip_decoded[7].t1 a_n1783_n1230# dvdd.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1056 comparator_0.vnn comparator_0.vpp avdd.t24 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1057 avdd.t184 comparator_0.vnn comparator_0.vnn avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1058 a_n20782_n2937# a_n20404_n10337# avss.t108 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1059 dvss.t376 a_10515_n2156# a_10874_n2222# dvss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1060 rc_osc_0.m rc_osc_0.in dvdd.t186 dvdd.t185 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X1061 a_n5214_n3990# a_n5639_n3946# dvss.t364 dvss.t363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1062 avdd.t270 avdd.t269 avdd.t270 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1063 a_n3102_n3990# a_n3527_n3946# dvss.t326 dvss.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1064 a_n990_n3990# a_n1415_n3946# dvss.t53 dvss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1065 vin_vunder.t30 avdd.t267 vin_vunder.t30 avdd.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1066 brout_filt.t18 sky130_fd_sc_hd__inv_4_0.Y dvss.t67 dvss.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1067 rstring_mux_0.vtrip1.t3 rstring_mux_0.otrip_decoded_avdd[1] vin_brout avss.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1068 rstring_mux_0.otrip_decoded_avdd[1] a_n6812_n1478# avdd.t154 avdd.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1069 rstring_mux_0.vtrip1.t7 rstring_mux_0.vtrip0.t5 avss.t257 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1070 dcomp.t3 sky130_fd_sc_hd__inv_4_3.Y dvdd.t297 dvdd.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1071 dvss.t250 a_10515_n1026# a_10874_n1026# dvss.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1072 a_n7326_n2256# a_n7751_n2212# dvss.t136 dvss.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1073 dvss.t595 a_n1683_n2876# a_n476_n3212# dvss.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1074 outb.t2 sky130_fd_sc_hd__inv_4_4.Y dvdd.t140 dvdd.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1075 a_10874_n2222# a_10515_n2156# dvss.t375 dvss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1076 avdd.t266 avdd.t263 avdd.t265 avdd.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=4
X1077 a_9145_n2212# a_8777_n1230# dvdd.t89 dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1078 dvss.t124 a_n6007_n2964# a_n5907_n2876# dvss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1079 a_n3649_n11914# rstring_mux_0.vtrip0.t0 avss.t156 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1080 avdd.t63 rstring_mux_0.ena_b rstring_mux_0.vtop.t3 avdd.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1081 sky130_fd_sc_hd__inv_4_3.Y vl dvdd.t69 dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1082 dvdd.t214 otrip_decoded[5].t1 a_n3895_n1230# dvdd.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1083 comparator_1.vt comparator_1.vn avss.t283 avss.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1084 a_10874_n1026# a_10515_n1026# dvss.t249 dvss.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1085 a_n7326_n3990# a_n7751_n3946# dvss.t5 dvss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1086 avdd.t262 avdd.t260 avdd.t261 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1087 a_697_n2212# a_329_n1230# dvdd.t225 dvdd.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1088 a_n8019_n2876# a_n8119_n2964# dvss.t207 dvss.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1089 dvdd.t170 vtrip_decoded[4].t1 a_4553_n2964# dvdd.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1090 avdd.t101 ibias_gen_0.vp.t12 comparator_0.ibias avdd.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1091 vunder.t18 sky130_fd_sc_hd__inv_4_1.Y dvss.t603 dvss.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1092 comparator_0.vnn comparator_0.vpp avdd.t23 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1093 avdd.t21 comparator_0.vpp comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1094 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1095 dcomp.t2 sky130_fd_sc_hd__inv_4_3.Y dvdd.t295 dvdd.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1096 a_1122_n3990# a_697_n3946# dvss.t442 dvss.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1097 vin_vunder.t46 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip1.t8 avss.t322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1098 ibg_200n comparator_0.ena a_n15479_n3901# avss.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X1099 avdd.t7 a_8877_n2876# a_9570_n3990# avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1100 a_4921_n3946# a_4553_n2964# dvdd.t97 dvdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1101 dcomp3v3uv comparator_0.n1 avss.t236 avss.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1102 avdd.t61 rstring_mux_0.ena_b rstring_mux_0.vtop.t2 avdd.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1103 avdd.t128 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1104 comparator_1.vpp vbg_1v2.t33 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1105 a_n16775_n2223# ibias_gen_0.ena_b ibias_gen_0.vstart.t0 avdd.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X1106 vin_vunder.t15 rstring_mux_0.vtrip_decoded_b_avdd[1] rstring_mux_0.vtrip1.t2 avdd.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1107 avdd.t510 ibias_gen_0.vp0.t12 ibias_gen_0.vn0.t16 avdd.t509 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1108 dvss.t316 a_2809_n3946# a_3234_n3990# dvss.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1109 comparator_1.vpp comparator_1.vnn avdd.t127 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1110 avdd.t589 comparator_1.n1 dcomp3v3 avdd.t588 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1111 dvss.t601 sky130_fd_sc_hd__inv_4_1.Y vunder.t17 dvss.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 dvdd.t200 otrip_decoded[3].t1 a_n6007_n1230# dvdd.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1113 dvss.t440 a_697_n3946# a_1122_n3990# dvss.t439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1114 ibias_gen_0.ve.t3 ibias_gen_0.vn0.t1 ibias_gen_0.vn0.t2 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1115 dvdd.t216 vtrip_decoded[6].t1 a_6665_n2964# dvdd.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1116 rstring_mux_0.vtrip3.t4 rstring_mux_0.otrip_decoded_b_avdd[3] vin_brout avdd.t500 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1117 a_2399_n11914# a_2021_n19314# avss.t157 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1118 a_n6673_n11914# a_n7051_n19314# avss.t104 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1119 avdd.t126 comparator_1.vnn comparator_1.vpp avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1120 vin_vunder.t37 rstring_mux_0.vtrip_decoded_avdd[0] rstring_mux_0.vtrip0.t8 avss.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1121 comparator_1.vnn comparator_1.vpp avdd.t459 avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1122 outb.t18 sky130_fd_sc_hd__inv_4_4.Y dvss.t391 dvss.t390 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1123 a_n7429_n11914# a_n7051_n19314# avss.t205 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1124 a_n10453_n11914# a_n10075_n19314# avss.t206 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1125 a_3234_n3990# a_2809_n3946# dvss.t314 dvss.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1126 dvss.t708 sky130_fd_sc_hd__inv_4_3.Y dcomp.t20 dvss.t707 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1127 rc_osc_0.in dvss.t479 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1128 avdd.t259 avdd.t257 avdd.t258 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1129 ibias_gen_0.vn0.t7 vbg_1v2.t34 ibias_gen_0.vstart.t2 avss.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1130 rc_osc_0.n.t4 rc_osc_0.m dvss.t657 dvss.t656 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1131 avdd.t458 comparator_1.vpp comparator_1.n0 avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1132 rstring_mux_0.vtrip_decoded_avdd[7] a_7972_n1478# avdd.t451 avdd.t450 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1133 dvdd.t202 otrip_decoded[1].t1 a_n8119_n1230# dvdd.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1134 dvss.t647 a_4921_n3946# a_5346_n3990# dvss.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1135 comparator_0.vnn avss.t392 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1136 a_n12731_9395# a_n13109_1995# avss.t303 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1137 avdd.t20 comparator_0.vpp comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1138 dvdd.t251 sky130_fd_sc_hd__inv_4_1.Y vunder.t9 dvdd.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1139 avdd.t256 avdd.t255 avdd.t256 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1140 dvdd.t182 outb_unbuf.t6 sky130_fd_sc_hd__inv_4_4.Y dvdd.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1141 schmitt_trigger_0.in.t11 dvss.t652 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1142 comparator_0.vpp vbg_1v2.t35 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1143 dvdd.t15 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t3 dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1144 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvdd.t227 dvdd.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1145 rstring_mux_0.vtrip6.t3 rstring_mux_0.otrip_decoded_avdd[6] vin_brout avss.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1146 avdd.t59 rstring_mux_0.ena_b rstring_mux_0.vtop.t1 avdd.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X1147 dvdd.t219 a_10874_n1026# a_10874_n2222# dvdd.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X1148 dvss.t381 a_429_n1142# a_1636_n1478# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1149 avdd.t497 a_n5907_n2876# a_n5214_n3990# avdd.t496 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1150 vin_brout avdd.t253 vin_brout avdd.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1151 rstring_mux_0.otrip_decoded_avdd[4] a_n2588_n3212# dvss.t535 dvss.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1152 a_5346_n3990# a_4921_n3946# dvss.t645 dvss.t644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1153 dvss.t232 a_10514_n2760# a_10514_n3890# dvss.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X1154 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.otrip_decoded_avdd[3] avdd.t582 avdd.t581 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1155 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip_decoded_avdd[0] avdd.t540 avdd.t539 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1156 dvdd.t184 rc_osc_0.in rc_osc_0.m dvdd.t183 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1157 dvss.t706 sky130_fd_sc_hd__inv_4_3.Y dcomp.t19 dvss.t705 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1158 ibias_gen_0.vn1.t6 ibias_gen_0.isrc_sel_b avss.t197 avss.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1159 avss.t34 avss.t33 avss.t34 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1160 dcomp.t1 sky130_fd_sc_hd__inv_4_3.Y dvdd.t293 dvdd.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 dvss.t247 a_10515_n1026# a_10874_n1026# dvss.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X1162 avdd.t542 comparator_0.ena rstring_mux_0.ena_b avdd.t541 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1163 osc_ck.t6 rc_osc_0.n.t13 dvdd.t223 dvdd.t222 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1164 vin_brout avss.t31 vin_brout avss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1165 outb.t1 sky130_fd_sc_hd__inv_4_4.Y dvdd.t138 dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1166 outb.t17 sky130_fd_sc_hd__inv_4_4.Y dvss.t389 dvss.t388 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1167 dvss.t346 a_7033_n3946# a_7458_n3990# dvss.t345 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1168 a_6179_n11914# a_5801_n19314# avss.t200 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1169 a_n13477_n11914# a_n13855_n19314# avss.t201 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1170 rstring_mux_0.otrip_decoded_avdd[1] a_n6812_n1478# dvss.t228 dvss.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1171 avdd.t252 avdd.t250 avdd.t251 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1172 vin_vunder.t24 avdd.t248 vin_vunder.t24 avdd.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1173 a_n8195_9395# a_n8573_1995# avss.t202 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1174 dvss.t102 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X sky130_fd_sc_hd__inv_4_1.A dvss.t101 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1175 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip_decoded_avdd[4] avdd.t409 avdd.t408 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1176 comparator_0.vm comparator_0.ena_b avss.t168 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1177 vin_vunder.t7 avss.t29 vin_brout avss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1178 sky130_fd_sc_hd__inv_4_3.Y vl dvdd.t67 dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1179 dvdd.t13 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t2 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1180 avdd.t19 comparator_0.vpp comparator_0.vpp avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1181 rstring_mux_0.otrip_decoded_avdd[7] a_n476_n1478# avdd.t173 avdd.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1182 comparator_0.vt vbg_1v2.t36 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1183 comparator_0.n0 comparator_0.vm avss.t337 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1184 avdd.t247 avdd.t245 avdd.t247 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1185 vin_brout avss.t27 vin_brout avss.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1186 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1187 avdd.t417 a_n8019_n2876# a_n7326_n3990# avdd.t416 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1188 brout_filt.t17 sky130_fd_sc_hd__inv_4_0.Y dvss.t65 dvss.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1189 a_2809_n3946# a_2441_n2964# dvss.t564 dvss.t563 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1190 avss.t26 avss.t23 avss.t25 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1191 dvss.t704 sky130_fd_sc_hd__inv_4_3.Y dcomp.t18 dvss.t703 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1192 dvss.t324 a_n3527_n3946# a_n3102_n3990# dvss.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1193 avss.t173 comparator_0.n0 comparator_0.n1 avss.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1194 vin_brout avss.t21 vin_brout avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1195 comparator_1.vnn vin_brout comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1196 avss.t124 comparator_0.vn comparator_0.vn avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1197 ibg_200n ibias_gen_0.ena_b a_n15529_n2223# avdd.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X1198 dvss.t150 a_9145_n3946# a_9570_n3990# dvss.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1199 a_887_n11914# a_1265_n19314# avss.t176 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1200 avdd.t427 comparator_0.n1 dcomp3v3uv avdd.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1201 comparator_1.vt avss.t393 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1202 a_n3102_n3990# a_n3527_n3946# dvss.t322 dvss.t321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1203 a_n10279_n23467# a_11121_n23089# dvss.t526 sky130_fd_pr__res_xhigh_po_1p41 l=105
X1204 dvdd.t11 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t1 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1205 rstring_mux_0.vtrip3.t1 rstring_mux_0.vtrip_decoded_avdd[3] vin_vunder.t10 avss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1206 dvss.t599 sky130_fd_sc_hd__inv_4_1.Y vunder.t16 dvss.t598 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1207 avdd.t244 avdd.t242 avdd.t243 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1208 dvss.t436 a_n3795_n2876# a_n2588_n3212# dvss.t435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1209 a_7033_n3946# a_6665_n2964# dvss.t583 dvss.t582 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1210 dvss.t362 a_n5639_n3946# a_n5214_n3990# dvss.t361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1211 schmitt_trigger_0.in.t12 dvss.t653 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1212 dvss.t280 a_4553_n2964# a_4653_n2876# dvss.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1213 rstring_mux_0.vtrip6.t8 rstring_mux_0.vtrip_decoded_avdd[6] vin_vunder.t35 avss.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1214 dvss.t310 otrip_decoded[6].t1 a_n1783_n2964# dvss.t309 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1215 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1216 comparator_0.vnn avss.t394 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1217 comparator_1.vt vin_brout comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1218 dvss.t454 outb_unbuf.t7 sky130_fd_sc_hd__inv_4_4.Y dvss.t453 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1219 comparator_0.vnn vin_vunder.t62 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1220 rstring_mux_0.vtrip1.t1 rstring_mux_0.vtrip_decoded_b_avdd[1] vin_vunder.t14 avdd.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1221 comparator_1.vpp comparator_1.vnn avdd.t124 avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1222 dcomp3v3uv comparator_0.n1 avss.t234 avss.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1223 comparator_0.vpp comparator_0.vnn avdd.t183 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1224 comparator_1.vpp vbg_1v2.t37 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1225 a_n5214_n3990# a_n5639_n3946# dvss.t360 dvss.t359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1226 schmitt_trigger_0.in.t13 dvss.t654 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1227 comparator_0.vpp vbg_1v2.t38 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1228 comparator_0.vnn avss.t395 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1229 avdd.t583 a_n1683_n1142# a_n476_n1478# avdd.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1230 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip_decoded_avdd[2] avss.t160 avss.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1231 comparator_0.vpp vbg_1v2.t39 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1232 dvdd.t136 sky130_fd_sc_hd__inv_4_4.Y outb.t0 dvdd.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1233 dvdd.t249 sky130_fd_sc_hd__inv_4_1.Y vunder.t1 dvdd.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1234 dvss.t537 a_n5907_n2876# a_n4700_n3212# dvss.t536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1235 vin_brout rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.vtrip3.t3 avdd.t499 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1236 a_4667_n11914# a_4289_n19314# avss.t177 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1237 dvss.t683 dvss.t681 rc_osc_0.n.t5 dvss.t682 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1238 a_1122_n3990# a_697_n3946# dvss.t438 dvss.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1239 a_9145_n3946# a_8777_n2964# dvss.t334 dvss.t333 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1240 a_n8941_n11914# a_n9319_n19314# avss.t203 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1241 a_n11965_n11914# a_n12343_n19314# avss.t204 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1242 comparator_1.n1 comparator_1.n0 avdd.t603 avdd.t602 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X1243 avdd.t241 avdd.t239 avdd.t241 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1244 avdd.t445 a_n990_n2256# a_n1683_n1142# avdd.t444 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1245 dvss.t3 a_n7751_n3946# a_n7326_n3990# dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1246 vin_vunder.t0 avss.t19 vin_vunder.t0 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1247 avdd.t238 avdd.t235 avdd.t237 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1248 avss.t226 comparator_1.vm comparator_1.vm avss.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1249 ibias_gen_0.vn0.t17 ibias_gen_0.vp0.t13 avdd.t512 avdd.t511 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1250 avss.t18 avss.t15 avss.t17 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X1251 a_4667_n11914# a_5045_n19314# avss.t221 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1252 comparator_0.vnn vin_vunder.t63 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1253 outb.t16 sky130_fd_sc_hd__inv_4_4.Y dvss.t387 dvss.t386 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1254 dvss.t226 otrip_decoded[4].t1 a_n3895_n2964# dvss.t225 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1255 schmitt_trigger_0.in.t14 dvss.t655 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1256 a_n12721_n11914# a_n12343_n19314# avss.t199 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1257 ibias_gen_0.vr.t1 avss.t13 ibias_gen_0.ve.t2 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1258 dvss.t702 sky130_fd_sc_hd__inv_4_3.Y dcomp.t17 dvss.t701 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1259 a_697_n3946# a_329_n2964# dvss.t294 dvss.t293 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1260 vin_brout avss.t11 vin_brout avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1261 ibias_gen_0.vp0.t0 avss.t9 ibias_gen_0.vn0.t0 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1262 rstring_mux_0.vtrip_decoded_avdd[4] a_5860_n3212# dvss.t560 dvss.t559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1263 ibias_gen_0.vn1.t8 avdd.t233 ibias_gen_0.vp1.t11 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1264 dvss.t518 schmitt_trigger_0.out.t15 sky130_fd_sc_hd__inv_4_0.Y dvss.t517 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1265 dcomp3v3uv comparator_0.n1 avdd.t425 avdd.t424 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1266 vin_brout avss.t7 vin_brout avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1267 comparator_1.vt vbg_1v2.t40 comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1268 avdd.t232 avdd.t230 avdd.t232 avdd.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X1269 avss.t6 avss.t4 avss.t6 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1270 dvdd.t247 sky130_fd_sc_hd__inv_4_1.Y vunder.t0 dvdd.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1271 dvss.t429 a_n8019_n2876# a_n6812_n3212# dvss.t428 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1272 avdd.t441 a_n3795_n2876# a_n3102_n3990# avdd.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1273 a_10514_n2760# dcomp3v3uv avdd.t49 avdd.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1274 avss.t3 avss.t1 avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1275 avdd.t229 avdd.t226 avdd.t228 avdd.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1276 dcomp3v3 comparator_1.n1 avdd.t587 avdd.t586 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1277 dcomp.t0 sky130_fd_sc_hd__inv_4_3.Y dvdd.t291 dvdd.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1278 dvdd.t9 sky130_fd_sc_hd__inv_4_0.Y brout_filt.t0 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1279 a_429_n2876# a_329_n2964# dvss.t292 dvss.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1280 a_3234_n3990# a_2809_n3946# dvss.t312 dvss.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1281 comparator_0.vt avss.t396 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1282 avdd.t182 comparator_0.vnn comparator_0.vm avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1283 a_10874_n1026# a_10874_n2222# dvdd.t204 dvdd.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X1284 dvss.t498 otrip_decoded[2].t1 a_n6007_n2964# dvss.t497 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1285 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.otrip_decoded_avdd[6] avss.t181 avss.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1286 ibias_gen_0.vstart.t1 vbg_1v2.t41 ibias_gen_0.vn0.t6 avss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1287 brout_filt.t16 sky130_fd_sc_hd__inv_4_0.Y dvss.t63 dvss.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1288 dvdd.t134 osc_ena.t3 rc_osc_0.in dvdd.t133 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X1289 comparator_0.vpp comparator_0.vnn avdd.t181 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1290 dvss.t700 sky130_fd_sc_hd__inv_4_3.Y dcomp.t16 dvss.t699 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1291 dvss.t643 a_4921_n3946# a_5346_n3990# dvss.t642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1292 schmitt_trigger_0.out.t3 schmitt_trigger_0.m.t17 dvss.t95 dvss.t94 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1293 comparator_1.vt avss.t397 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1294 dvss.t173 a_429_n2876# a_1636_n3212# dvss.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
R0 avss.n68 avss.n67 2.18688e+07
R1 avss.n370 avss.n369 188352
R2 avss.n671 avss.n635 160432
R3 avss.n635 avss.n634 110760
R4 avss.n66 avss.n50 100279
R5 avss.n797 avss.n50 100279
R6 avss.n66 avss.n51 100279
R7 avss.n797 avss.n51 100279
R8 avss.n369 avss.n368 92956.3
R9 avss.n308 avss.n69 68021.9
R10 avss.n781 avss.n363 64733.3
R11 avss.n369 avss.t174 48414.6
R12 avss.n660 avss.n360 45524.4
R13 avss.n660 avss.n361 45524.4
R14 avss.n783 avss.n360 45524.4
R15 avss.n783 avss.n361 45524.4
R16 avss.n568 avss.n563 45524.4
R17 avss.n632 avss.n563 45524.4
R18 avss.n568 avss.n565 45524.4
R19 avss.n632 avss.n565 45524.4
R20 avss.n308 avss.n307 45183
R21 avss.n880 avss.n8 37415.6
R22 avss.n781 avss.n780 29160.7
R23 avss.n635 avss.t360 29031.2
R24 avss.n800 avss.n47 21059.4
R25 avss.n800 avss.n48 21059.4
R26 avss.n802 avss.n47 21059.4
R27 avss.n802 avss.n48 21059.4
R28 avss.n766 avss.n372 18174.6
R29 avss.n773 avss.n372 18174.6
R30 avss.n773 avss.n371 18174.6
R31 avss.n766 avss.n371 18174.6
R32 avss.n617 avss.n553 18174.6
R33 avss.n589 avss.n553 18174.6
R34 avss.n617 avss.n616 18174.6
R35 avss.n616 avss.n589 18174.6
R36 avss.n344 avss.n63 16300.9
R37 avss.n340 avss.n63 16300.9
R38 avss.n344 avss.n65 16300.9
R39 avss.n340 avss.n65 16300.9
R40 avss.n672 avss.n671 13864
R41 avss.n117 avss.n69 12588.9
R42 avss.n669 avss.n637 12517.1
R43 avss.n663 avss.n637 12517.1
R44 avss.n663 avss.n636 12517.1
R45 avss.n669 avss.n636 12517.1
R46 avss.n443 avss.n439 7742.83
R47 avss.n445 avss.n439 7742.83
R48 avss.n444 avss.n443 7742.83
R49 avss.n445 avss.n444 7742.83
R50 avss.n650 avss.n19 7610.36
R51 avss.n650 avss.n20 7610.36
R52 avss.n857 avss.n20 7610.36
R53 avss.n857 avss.n19 7610.36
R54 avss.n54 avss.n52 6515.58
R55 avss.n796 avss.n52 6515.58
R56 avss.n795 avss.n54 6515.58
R57 avss.n796 avss.n795 6515.58
R58 avss.n860 avss.n12 5644.38
R59 avss.n860 avss.n13 5644.38
R60 avss.n871 avss.n13 5644.38
R61 avss.n871 avss.n12 5644.38
R62 avss.n69 avss.n68 4523.98
R63 avss.n442 avss.n437 4175.68
R64 avss.n446 avss.n437 4175.68
R65 avss.n442 avss.n438 4175.68
R66 avss.n446 avss.n438 4175.68
R67 avss.n760 avss.n379 4139.43
R68 avss.n756 avss.n379 4139.43
R69 avss.n760 avss.n380 4139.43
R70 avss.n756 avss.n380 4139.43
R71 avss.n621 avss.n582 4139.43
R72 avss.n587 avss.n582 4139.43
R73 avss.n587 avss.n583 4139.43
R74 avss.n621 avss.n583 4139.43
R75 avss.n561 avss.n557 3978.07
R76 avss.n561 avss.n558 3978.07
R77 avss.n675 avss.n558 3978.07
R78 avss.n675 avss.n557 3978.07
R79 avss.n779 avss.n365 3978.07
R80 avss.n775 avss.n365 3978.07
R81 avss.n775 avss.n364 3978.07
R82 avss.n779 avss.n364 3978.07
R83 avss.t229 avss.t40 3966.94
R84 avss.t227 avss.t229 3966.94
R85 avss.t225 avss.t231 3966.94
R86 avss.t231 avss.t61 3966.94
R87 avss.n874 avss.n9 3902.33
R88 avss.n874 avss.n10 3902.33
R89 avss.n878 avss.n10 3902.33
R90 avss.n878 avss.n9 3902.33
R91 avss.n671 avss.n670 3318.88
R92 avss.n322 avss.n321 2998.14
R93 avss.n784 avss.n359 2957.93
R94 avss.n631 avss.n566 2957.93
R95 avss.n630 avss.n569 2957.93
R96 avss.n631 avss.n630 2957.93
R97 avss.n626 avss.n569 2940.24
R98 avss.n659 avss.n359 2935.34
R99 avss.n129 avss.n128 2905.02
R100 avss.n141 avss.n140 2905.02
R101 avss.n153 avss.n152 2905.02
R102 avss.n165 avss.n164 2905.02
R103 avss.n177 avss.n176 2905.02
R104 avss.n189 avss.n188 2905.02
R105 avss.n201 avss.n200 2905.02
R106 avss.n213 avss.n212 2905.02
R107 avss.n225 avss.n224 2905.02
R108 avss.n237 avss.n236 2905.02
R109 avss.n249 avss.n248 2905.02
R110 avss.n261 avss.n260 2905.02
R111 avss.n273 avss.n272 2905.02
R112 avss.n285 avss.n284 2905.02
R113 avss.n297 avss.n296 2905.02
R114 avss.n882 avss.n881 2538.7
R115 avss.t356 avss.n582 2436.62
R116 avss.n583 avss.t360 2436.62
R117 avss.n379 avss.t241 2436.62
R118 avss.n803 avss.n45 2366.87
R119 avss.n803 avss.n44 2366.87
R120 avss.n799 avss.n44 2344.28
R121 avss.n799 avss.n45 2344.28
R122 avss.n618 avss.t40 2304.08
R123 avss.t61 avss.n562 2304.08
R124 avss.n489 avss.n473 2087.09
R125 avss.n514 avss.n463 2084.98
R126 avss.n614 avss.n552 2054.02
R127 avss.n679 avss.n552 2054.02
R128 avss.n772 avss.n373 2054.02
R129 avss.n767 avss.n373 2054.02
R130 avss.n507 avss.n505 2039.85
R131 avss.n531 avss.n530 2039.84
R132 avss.n615 avss.t227 1983.47
R133 avss.n615 avss.t225 1983.47
R134 avss.n679 avss.n678 1894.78
R135 avss.n614 avss.n590 1894.78
R136 avss.n769 avss.n767 1894.78
R137 avss.n772 avss.n771 1894.78
R138 avss.n339 avss.n338 1813.84
R139 avss.n884 avss.n6 1735.47
R140 avss.n885 avss.n6 1735.47
R141 avss.n885 avss.n5 1735.47
R142 avss.n884 avss.n5 1735.47
R143 avss.t235 avss.n49 1637.21
R144 avss.n346 avss.n62 1602.64
R145 avss.n653 avss.n652 1487.81
R146 avss.n652 avss.n357 1487.81
R147 avss.n659 avss.n653 1439.24
R148 avss.n784 avss.n357 1439.24
R149 avss.n664 avss.n649 1435.48
R150 avss.n664 avss.n648 1435.48
R151 avss.n321 avss.n320 1414.29
R152 avss.t293 avss.t302 1389.88
R153 avss.n668 avss.n639 1385.79
R154 avss.n668 avss.n638 1385.79
R155 avss.n620 avss.t344 1301
R156 avss.n620 avss.t348 1301
R157 avss.n761 avss.t237 1301
R158 avss.t247 avss.n761 1301
R159 avss.n780 avss.t302 1143.92
R160 avss.t348 avss.t354 1081.77
R161 avss.t241 avss.t233 1081.77
R162 avss.t346 avss.t356 1081.77
R163 avss.t350 avss.t346 1081.77
R164 avss.t352 avss.t350 1081.77
R165 avss.t344 avss.t352 1081.77
R166 avss.t354 avss.t342 1081.77
R167 avss.t342 avss.t358 1081.77
R168 avss.t233 avss.t245 1081.77
R169 avss.t245 avss.t243 1081.77
R170 avss.n441 avss.n434 976.942
R171 avss.n441 avss.n440 976.942
R172 avss.n448 avss.n447 976.188
R173 avss.n447 avss.n436 974.683
R174 avss.t172 avss.n49 964.784
R175 avss.n321 avss.n308 939.895
R176 avss.n588 avss.t344 925.769
R177 avss.t348 avss.n588 925.769
R178 avss.n619 avss.t360 887.293
R179 avss.n856 avss.n21 874.542
R180 avss.n22 avss.n21 874.542
R181 avss.n128 avss.n115 815.444
R182 avss.n140 avss.n112 815.444
R183 avss.n152 avss.n109 815.444
R184 avss.n164 avss.n106 815.444
R185 avss.n176 avss.n103 815.444
R186 avss.n188 avss.n100 815.444
R187 avss.n200 avss.n97 815.444
R188 avss.n212 avss.n94 815.444
R189 avss.n224 avss.n91 815.444
R190 avss.n236 avss.n88 815.444
R191 avss.n248 avss.n85 815.444
R192 avss.n260 avss.n82 815.444
R193 avss.n272 avss.n79 815.444
R194 avss.n284 avss.n76 815.444
R195 avss.n296 avss.n73 815.444
R196 avss.n307 avss.n70 815.444
R197 avss.n59 avss.n58 796.612
R198 avss.n64 avss.n58 782.683
R199 avss.n312 avss.n309 769.572
R200 avss.n854 avss.n853 765.741
R201 avss.n855 avss.n854 765.741
R202 avss.n56 avss.n55 759.718
R203 avss.n117 avss.t307 755.986
R204 avss.n129 avss.t275 755.986
R205 avss.n141 avss.t110 755.986
R206 avss.n153 avss.t217 755.986
R207 avss.n165 avss.t132 755.986
R208 avss.n177 avss.t159 755.986
R209 avss.n189 avss.t323 755.986
R210 avss.n201 avss.t290 755.986
R211 avss.n213 avss.t363 755.986
R212 avss.n225 avss.t180 755.986
R213 avss.n237 avss.t153 755.986
R214 avss.n249 avss.t329 755.986
R215 avss.n261 avss.t332 755.986
R216 avss.n273 avss.t137 755.986
R217 avss.n285 avss.t189 755.986
R218 avss.n297 avss.t277 755.986
R219 avss.t297 avss.t295 731.963
R220 avss.t265 avss.t269 731.963
R221 avss.t269 avss.n673 684.673
R222 avss.n674 avss.t295 668.225
R223 avss.n870 avss.n14 649.788
R224 avss.n861 avss.n14 649.788
R225 avss.n782 avss.n781 627.813
R226 avss.n506 avss.t43 625.516
R227 avss.n513 avss.t43 625.516
R228 avss.t43 avss.n457 614.321
R229 avss.n524 avss.t43 614.321
R230 avss.n634 avss.t297 602.431
R231 avss.n57 avss.n56 598.966
R232 avss.t43 avss.n496 598.606
R233 avss.n497 avss.t43 598.606
R234 avss.n482 avss.t43 588.343
R235 avss.n480 avss.t43 588.343
R236 avss.n319 avss.n318 585
R237 avss.n320 avss.n319 585
R238 avss.n311 avss.n310 585
R239 avss.n503 avss.n502 585
R240 avss.n501 avss.n470 585
R241 avss.n470 avss.n469 585
R242 avss.n500 avss.n499 585
R243 avss.n499 avss.n498 585
R244 avss.n472 avss.n471 585
R245 avss.n497 avss.n472 585
R246 avss.n495 avss.n494 585
R247 avss.n496 avss.n495 585
R248 avss.n493 avss.n474 585
R249 avss.n474 avss.n473 585
R250 avss.n492 avss.n491 585
R251 avss.n476 avss.n475 585
R252 avss.n518 avss.n517 585
R253 avss.n515 avss.n465 585
R254 avss.n515 avss.n514 585
R255 avss.n512 avss.n511 585
R256 avss.n513 avss.n512 585
R257 avss.n510 avss.n466 585
R258 avss.n506 avss.n466 585
R259 avss.n509 avss.n508 585
R260 avss.n508 avss.n507 585
R261 avss.n468 avss.n467 585
R262 avss.n519 avss.n464 585
R263 avss.n521 avss.n520 585
R264 avss.n522 avss.n521 585
R265 avss.n462 avss.n461 585
R266 avss.n523 avss.n462 585
R267 avss.n526 avss.n525 585
R268 avss.n525 avss.n524 585
R269 avss.n527 avss.n459 585
R270 avss.n459 avss.n457 585
R271 avss.n529 avss.n528 585
R272 avss.n530 avss.n529 585
R273 avss.n460 avss.n458 585
R274 avss.n454 avss.n452 585
R275 avss.n487 avss.n486 585
R276 avss.n488 avss.n487 585
R277 avss.n485 avss.n478 585
R278 avss.n478 avss.n477 585
R279 avss.n484 avss.n483 585
R280 avss.n483 avss.n482 585
R281 avss.n481 avss.n479 585
R282 avss.n481 avss.n480 585
R283 avss.n453 avss.n451 585
R284 avss.n455 avss.n453 585
R285 avss.n534 avss.n533 585
R286 avss.n533 avss.n532 585
R287 avss.n119 avss.n118 585
R288 avss.n118 avss.n117 585
R289 avss.n120 avss.n116 585
R290 avss.n116 avss.n115 585
R291 avss.n127 avss.n126 585
R292 avss.n128 avss.n127 585
R293 avss.n131 avss.n130 585
R294 avss.n130 avss.n129 585
R295 avss.n114 avss.n113 585
R296 avss.n113 avss.n112 585
R297 avss.n139 avss.n138 585
R298 avss.n140 avss.n139 585
R299 avss.n143 avss.n142 585
R300 avss.n142 avss.n141 585
R301 avss.n111 avss.n110 585
R302 avss.n110 avss.n109 585
R303 avss.n151 avss.n150 585
R304 avss.n152 avss.n151 585
R305 avss.n155 avss.n154 585
R306 avss.n154 avss.n153 585
R307 avss.n108 avss.n107 585
R308 avss.n107 avss.n106 585
R309 avss.n163 avss.n162 585
R310 avss.n164 avss.n163 585
R311 avss.n167 avss.n166 585
R312 avss.n166 avss.n165 585
R313 avss.n105 avss.n104 585
R314 avss.n104 avss.n103 585
R315 avss.n175 avss.n174 585
R316 avss.n176 avss.n175 585
R317 avss.n179 avss.n178 585
R318 avss.n178 avss.n177 585
R319 avss.n102 avss.n101 585
R320 avss.n101 avss.n100 585
R321 avss.n187 avss.n186 585
R322 avss.n188 avss.n187 585
R323 avss.n191 avss.n190 585
R324 avss.n190 avss.n189 585
R325 avss.n99 avss.n98 585
R326 avss.n98 avss.n97 585
R327 avss.n199 avss.n198 585
R328 avss.n200 avss.n199 585
R329 avss.n203 avss.n202 585
R330 avss.n202 avss.n201 585
R331 avss.n96 avss.n95 585
R332 avss.n95 avss.n94 585
R333 avss.n211 avss.n210 585
R334 avss.n212 avss.n211 585
R335 avss.n215 avss.n214 585
R336 avss.n214 avss.n213 585
R337 avss.n93 avss.n92 585
R338 avss.n92 avss.n91 585
R339 avss.n223 avss.n222 585
R340 avss.n224 avss.n223 585
R341 avss.n227 avss.n226 585
R342 avss.n226 avss.n225 585
R343 avss.n90 avss.n89 585
R344 avss.n89 avss.n88 585
R345 avss.n235 avss.n234 585
R346 avss.n236 avss.n235 585
R347 avss.n239 avss.n238 585
R348 avss.n238 avss.n237 585
R349 avss.n87 avss.n86 585
R350 avss.n86 avss.n85 585
R351 avss.n247 avss.n246 585
R352 avss.n248 avss.n247 585
R353 avss.n251 avss.n250 585
R354 avss.n250 avss.n249 585
R355 avss.n84 avss.n83 585
R356 avss.n83 avss.n82 585
R357 avss.n259 avss.n258 585
R358 avss.n260 avss.n259 585
R359 avss.n263 avss.n262 585
R360 avss.n262 avss.n261 585
R361 avss.n81 avss.n80 585
R362 avss.n80 avss.n79 585
R363 avss.n271 avss.n270 585
R364 avss.n272 avss.n271 585
R365 avss.n275 avss.n274 585
R366 avss.n274 avss.n273 585
R367 avss.n78 avss.n77 585
R368 avss.n77 avss.n76 585
R369 avss.n283 avss.n282 585
R370 avss.n284 avss.n283 585
R371 avss.n287 avss.n286 585
R372 avss.n286 avss.n285 585
R373 avss.n75 avss.n74 585
R374 avss.n74 avss.n73 585
R375 avss.n295 avss.n294 585
R376 avss.n296 avss.n295 585
R377 avss.n299 avss.n298 585
R378 avss.n298 avss.n297 585
R379 avss.n72 avss.n71 585
R380 avss.n71 avss.n70 585
R381 avss.n306 avss.n305 585
R382 avss.n307 avss.n306 585
R383 avss.n862 avss.n15 540.989
R384 avss.n869 avss.n15 540.989
R385 avss.n319 avss.n310 539.294
R386 avss.n298 avss.n71 539.294
R387 avss.n306 avss.n71 539.294
R388 avss.n286 avss.n74 539.294
R389 avss.n295 avss.n74 539.294
R390 avss.n274 avss.n77 539.294
R391 avss.n283 avss.n77 539.294
R392 avss.n262 avss.n80 539.294
R393 avss.n271 avss.n80 539.294
R394 avss.n250 avss.n83 539.294
R395 avss.n259 avss.n83 539.294
R396 avss.n238 avss.n86 539.294
R397 avss.n247 avss.n86 539.294
R398 avss.n226 avss.n89 539.294
R399 avss.n235 avss.n89 539.294
R400 avss.n214 avss.n92 539.294
R401 avss.n223 avss.n92 539.294
R402 avss.n202 avss.n95 539.294
R403 avss.n211 avss.n95 539.294
R404 avss.n190 avss.n98 539.294
R405 avss.n199 avss.n98 539.294
R406 avss.n178 avss.n101 539.294
R407 avss.n187 avss.n101 539.294
R408 avss.n166 avss.n104 539.294
R409 avss.n175 avss.n104 539.294
R410 avss.n154 avss.n107 539.294
R411 avss.n163 avss.n107 539.294
R412 avss.n142 avss.n110 539.294
R413 avss.n151 avss.n110 539.294
R414 avss.n130 avss.n113 539.294
R415 avss.n139 avss.n113 539.294
R416 avss.n118 avss.n116 539.294
R417 avss.n127 avss.n116 539.294
R418 avss.n321 avss.t300 492.382
R419 avss.n378 avss.t293 488.039
R420 avss.n586 avss.n581 477.741
R421 avss.n622 avss.n581 477.741
R422 avss.n758 avss.n757 477.741
R423 avss.n759 avss.n758 477.741
R424 avss.t267 avss.n672 474.954
R425 avss.n676 avss.n556 459.295
R426 avss.n560 avss.n556 459.295
R427 avss.n560 avss.n559 459.295
R428 avss.n778 avss.n366 459.295
R429 avss.n778 avss.n777 459.295
R430 avss.n777 avss.n776 459.295
R431 avss.n483 avss.n481 456.416
R432 avss.n525 avss.n459 456.416
R433 avss.n512 avss.n466 456.416
R434 avss.n495 avss.n472 456.416
R435 avss.n877 avss.n11 425.264
R436 avss.n875 avss.n11 420.43
R437 avss.n876 avss.n875 420.43
R438 avss.n877 avss.n876 420.43
R439 avss.n623 avss.n580 401.812
R440 avss.n585 avss.n580 401.812
R441 avss.n382 avss.n381 401.812
R442 avss.n755 avss.n382 401.812
R443 avss.n25 avss.t9 392.769
R444 avss.n24 avss.t81 392.692
R445 avss.n23 avss.t53 392.664
R446 avss.n61 avss.t19 384.515
R447 avss.n323 avss.t77 384.515
R448 avss.n325 avss.t73 384.515
R449 avss.n326 avss.t79 384.515
R450 avss.n327 avss.t75 384.515
R451 avss.n328 avss.t51 384.515
R452 avss.n329 avss.t29 384.515
R453 avss.n336 avss.t7 384.515
R454 avss.n334 avss.t31 384.515
R455 avss.n333 avss.t11 384.515
R456 avss.n332 avss.t64 384.515
R457 avss.n331 avss.t27 384.515
R458 avss.n330 avss.t55 384.515
R459 avss.n324 avss.t83 384.454
R460 avss.n335 avss.t21 384.454
R461 avss.n661 avss.t115 382.757
R462 avss.n507 avss.n506 363.548
R463 avss.n514 avss.n513 363.548
R464 avss.n530 avss.n457 357.041
R465 avss.n524 avss.n523 357.041
R466 avss.n523 avss.n522 357.041
R467 avss.n522 avss.n463 357.041
R468 avss.n496 avss.n473 347.908
R469 avss.n498 avss.n497 347.908
R470 avss.n498 avss.n469 347.908
R471 avss.n505 avss.n469 347.908
R472 avss.n489 avss.n488 341.943
R473 avss.n488 avss.n477 341.943
R474 avss.n482 avss.n477 341.943
R475 avss.n480 avss.n455 341.943
R476 avss.n532 avss.n455 341.943
R477 avss.n532 avss.n531 341.943
R478 avss.n619 avss.n618 340.805
R479 avss.n363 avss.t108 338.375
R480 avss.n419 avss.n406 333.334
R481 avss.n414 avss.n413 333.334
R482 avss.n429 avss.n404 333.334
R483 avss.t120 avss.n7 323.332
R484 avss.t120 avss.n882 323.332
R485 avss.n677 avss.n555 318.495
R486 avss.n768 avss.n367 318.495
R487 avss.n321 avss.n7 301.202
R488 avss.n516 avss.n463 283.521
R489 avss.n505 avss.n504 283.521
R490 avss.n339 avss.n55 274.072
R491 avss.n345 avss.n59 270.683
R492 avss.n670 avss.t14 262.885
R493 avss.n662 avss.t14 262.885
R494 avss.n490 avss.n489 262.719
R495 avss.n531 avss.n456 262.719
R496 avss.n782 avss.t16 239.365
R497 avss.n346 avss.n345 238.306
R498 avss.n673 avss.n562 227.298
R499 avss.t88 avss.n11 209.756
R500 avss.n876 avss.t88 209.756
R501 avss.n64 avss.n57 208.189
R502 avss.n883 avss.n4 202.918
R503 avss.n886 avss.n4 202.918
R504 avss.n320 avss.n309 200.215
R505 avss.t358 avss.n619 194.476
R506 avss.n883 avss.n3 193.918
R507 avss.n651 avss.t16 188.975
R508 avss.n887 avss.n886 186.73
R509 avss.t105 avss.t251 185.605
R510 avss.t251 avss.t335 185.605
R511 avss.t335 avss.t123 185.605
R512 avss.t123 avss.t104 185.605
R513 avss.t104 avss.t205 185.605
R514 avss.t205 avss.t122 185.605
R515 avss.t122 avss.t271 185.605
R516 avss.t271 avss.t254 185.605
R517 avss.n424 avss.n423 185
R518 avss.n425 avss.n411 185
R519 avss.n417 avss.n416 185
R520 avss.n418 avss.n406 185
R521 avss.t42 avss.n406 185
R522 avss.n420 avss.n419 185
R523 avss.n422 avss.n421 185
R524 avss.n413 avss.n412 185
R525 avss.n415 avss.n414 185
R526 avss.n405 avss.n403 185
R527 avss.n430 avss.n429 185
R528 avss.n429 avss.t42 185
R529 avss.n404 avss.n402 185
R530 avss.n427 avss.n426 185
R531 avss.n310 avss.n309 184.572
R532 avss.t224 avss.t312 160.339
R533 avss.t139 avss.t224 160.339
R534 avss.t220 avss.t139 160.339
R535 avss.t101 avss.t220 160.339
R536 avss.t255 avss.t253 160.339
R537 avss.t253 avss.t116 160.339
R538 avss.t116 avss.t193 160.339
R539 avss.t193 avss.t191 160.339
R540 avss.t191 avss.t200 160.339
R541 avss.t200 avss.t222 160.339
R542 avss.t222 avss.t194 160.339
R543 avss.t194 avss.t221 160.339
R544 avss.t221 avss.t177 160.339
R545 avss.t177 avss.t109 160.339
R546 avss.n678 avss.n554 159.248
R547 avss.n590 avss.n554 159.248
R548 avss.n770 avss.n769 159.248
R549 avss.n771 avss.n770 159.248
R550 avss.n68 avss.t101 157.37
R551 avss.n316 avss.t301 149.067
R552 avss.n302 avss.t278 149.067
R553 avss.n291 avss.t190 149.067
R554 avss.n279 avss.t138 149.067
R555 avss.n267 avss.t333 149.067
R556 avss.n255 avss.t330 149.067
R557 avss.n243 avss.t154 149.067
R558 avss.n231 avss.t181 149.067
R559 avss.n219 avss.t364 149.067
R560 avss.n207 avss.t291 149.067
R561 avss.n195 avss.t324 149.067
R562 avss.n183 avss.t160 149.067
R563 avss.n171 avss.t133 149.067
R564 avss.n159 avss.t218 149.067
R565 avss.n147 avss.t111 149.067
R566 avss.n135 avss.t276 149.067
R567 avss.n123 avss.t308 149.067
R568 avss.n341 avss.t213 142.101
R569 avss.n322 avss.t105 132.919
R570 avss.n487 avss.n478 132.635
R571 avss.n483 avss.n478 132.635
R572 avss.n481 avss.n453 132.635
R573 avss.n533 avss.n453 132.635
R574 avss.n529 avss.n458 132.635
R575 avss.n529 avss.n459 132.635
R576 avss.n525 avss.n462 132.635
R577 avss.n521 avss.n462 132.635
R578 avss.n521 avss.n464 132.635
R579 avss.n508 avss.n468 132.635
R580 avss.n508 avss.n466 132.635
R581 avss.n515 avss.n512 132.635
R582 avss.n517 avss.n515 132.635
R583 avss.n491 avss.n474 132.635
R584 avss.n495 avss.n474 132.635
R585 avss.n499 avss.n472 132.635
R586 avss.n499 avss.n470 132.635
R587 avss.n503 avss.n470 132.635
R588 avss.t321 avss.t202 132.379
R589 avss.t202 avss.t100 132.379
R590 avss.t100 avss.t150 132.379
R591 avss.t150 avss.t259 132.379
R592 avss.t195 avss.t264 132.379
R593 avss.t287 avss.t195 132.379
R594 avss.t309 avss.t287 132.379
R595 avss.t106 avss.t309 132.379
R596 avss.t117 avss.t140 132.379
R597 avss.t140 avss.t107 132.379
R598 avss.t107 avss.t303 132.379
R599 avss.t303 avss.t184 132.379
R600 avss.t184 avss.t223 132.379
R601 avss.t223 avss.t207 132.379
R602 avss.t207 avss.t118 132.379
R603 avss.t118 avss.t263 132.379
R604 avss.t263 avss.t311 132.379
R605 avss.n635 avss.n633 129.577
R606 avss.t143 avss.n49 118.332
R607 avss.t256 avss.t203 118.26
R608 avss.t203 avss.t98 118.26
R609 avss.t98 avss.t211 118.26
R610 avss.t211 avss.t206 118.26
R611 avss.t206 avss.t210 118.26
R612 avss.n582 avss.n580 117.001
R613 avss.n583 avss.n581 117.001
R614 avss.n557 avss.n556 117.001
R615 avss.n634 avss.n557 117.001
R616 avss.n559 avss.n558 117.001
R617 avss.n672 avss.n558 117.001
R618 avss.n779 avss.n778 117.001
R619 avss.n780 avss.n779 117.001
R620 avss.n758 avss.n380 117.001
R621 avss.n380 avss.n370 117.001
R622 avss.n776 avss.n775 117.001
R623 avss.n775 avss.n774 117.001
R624 avss.n382 avss.n379 117.001
R625 avss.n884 avss.n883 117.001
R626 avss.t120 avss.n884 117.001
R627 avss.n886 avss.n885 117.001
R628 avss.n885 avss.t120 117.001
R629 avss.n416 avss.n406 113.334
R630 avss.n429 avss.n405 113.334
R631 avss.n662 avss.n661 111.906
R632 avss.t210 avss.t167 110.1
R633 avss.t312 avss.n67 107.742
R634 avss.n559 avss.n555 99.0123
R635 avss.n776 avss.n367 99.0123
R636 avss.n5 avss.n3 97.5005
R637 avss.n7 avss.n5 97.5005
R638 avss.n6 avss.n4 97.5005
R639 avss.n882 avss.n6 97.5005
R640 avss.t212 avss.t314 96.6926
R641 avss.n343 avss.t305 94.5922
R642 avss.n568 avss.t321 93.9962
R643 avss.t165 avss.t201 91.065
R644 avss.n633 avss.t311 88.9531
R645 avss.n571 avss.t357 88.2028
R646 avss.n575 avss.t361 88.2028
R647 avss.n714 avss.t169 88.2028
R648 avss.n384 avss.t242 88.2028
R649 avss.n388 avss.t175 88.2028
R650 avss.n683 avss.t268 88.2028
R651 avss.n716 avss.t294 87.8727
R652 avss.n685 avss.t296 87.8727
R653 avss.n411 avss.n409 87.6787
R654 avss.n423 avss.n409 87.6787
R655 avss.n715 avss.t171 87.5075
R656 avss.n714 avss.t168 87.5075
R657 avss.n684 avss.t266 87.5075
R658 avss.n683 avss.t270 87.5075
R659 avss.n856 avss.n855 86.2123
R660 avss.n853 avss.n22 86.2123
R661 avss.n870 avss.n869 86.2123
R662 avss.n862 avss.n861 86.2123
R663 avss.n888 avss.t121 85.1191
R664 avss.t167 avss.n880 84.4142
R665 avss.n688 avss.t72 82.9912
R666 avss.n540 avss.t63 82.9912
R667 avss.n596 avss.t47 82.9912
R668 avss.t41 avss.n607 82.9912
R669 avss.t3 avss.n747 82.9912
R670 avss.t45 avss.n744 82.9912
R671 avss.n719 avss.t87 82.9912
R672 avss.n706 avss.t26 82.9912
R673 avss.n678 avss.n677 82.824
R674 avss.n590 avss.n555 82.824
R675 avss.n769 avss.n768 82.824
R676 avss.n771 avss.n367 82.824
R677 avss.t179 avss.t163 81.8562
R678 avss.t264 avss.n8 79.8477
R679 avss.t42 avss.n407 77.7851
R680 avss.t42 avss.n408 77.7851
R681 avss.t279 avss.t258 76.3526
R682 avss.t306 avss.t20 75.5042
R683 avss.t274 avss.t273 75.5042
R684 avss.t78 avss.t113 75.5042
R685 avss.t112 avss.t84 75.5042
R686 avss.t216 avss.t219 75.5042
R687 avss.t74 avss.t134 75.5042
R688 avss.t134 avss.t131 75.5042
R689 avss.t80 avss.t161 75.5042
R690 avss.t162 avss.t76 75.5042
R691 avss.t322 avss.t325 75.5042
R692 avss.t52 avss.t288 75.5042
R693 avss.t289 avss.t30 75.5042
R694 avss.t362 avss.t365 75.5042
R695 avss.t8 avss.t183 75.5042
R696 avss.t182 avss.t22 75.5042
R697 avss.t22 avss.t152 75.5042
R698 avss.t155 avss.t32 75.5042
R699 avss.t328 avss.t327 75.5042
R700 avss.t12 avss.t331 75.5042
R701 avss.t334 avss.t65 75.5042
R702 avss.t28 avss.t188 75.5042
R703 avss.t187 avss.t56 75.5042
R704 avss.t280 avss.t279 75.5042
R705 avss.t208 avss.t155 73.8075
R706 avss.n881 avss.t254 73.162
R707 avss.t0 avss.t80 72.9591
R708 avss.n881 avss.t256 71.6444
R709 avss.n573 avss.n572 70.9775
R710 avss.n571 avss.n570 70.9775
R711 avss.n577 avss.n576 70.9775
R712 avss.n575 avss.n574 70.9775
R713 avss.n386 avss.n385 70.9775
R714 avss.n384 avss.n383 70.9775
R715 avss.n390 avss.n389 70.9775
R716 avss.n388 avss.n387 70.9775
R717 avss.n546 avss.n545 70.9612
R718 avss.n544 avss.n543 70.9612
R719 avss.n550 avss.n549 70.9612
R720 avss.n612 avss.n611 70.9612
R721 avss.n595 avss.n592 70.9612
R722 avss.n609 avss.n608 70.9612
R723 avss.n712 avss.n711 70.9612
R724 avss.n710 avss.n709 70.9612
R725 avss.n396 avss.n395 70.9612
R726 avss.n394 avss.n393 70.9612
R727 avss.n749 avss.n748 70.9612
R728 avss.n746 avss.n745 70.9612
R729 avss.t42 avss.n410 70.8113
R730 avss.t42 avss.n428 70.8113
R731 avss.t317 avss.t252 70.601
R732 avss.n423 avss.n422 70.0005
R733 avss.n427 avss.n411 70.0005
R734 avss.t219 avss.t310 68.7174
R735 avss.t282 avss.t114 67.9453
R736 avss.t281 avss.t282 67.9453
R737 avss.t115 avss.t281 67.9453
R738 avss.t183 avss.t192 67.869
R739 avss.t56 avss.t178 67.0206
R740 avss.n564 avss.t106 66.1896
R741 avss.n564 avss.t117 66.1896
R742 avss.t336 avss.t328 64.4756
R743 avss.t247 avss.t239 63.8987
R744 avss.n674 avss.t265 63.7388
R745 avss.t176 avss.t162 63.6272
R746 avss.n378 avss.t237 63.1818
R747 avss.n363 avss.n362 61.8334
R748 avss.t151 avss.t196 61.3923
R749 avss.n873 avss.t5 61.1365
R750 avss.n879 avss.t204 60.3691
R751 avss.n458 avss.n456 59.5655
R752 avss.n491 avss.n490 59.5655
R753 avss.n490 avss.n476 59.5655
R754 avss.n456 avss.n454 59.5655
R755 avss.t307 avss.n115 59.46
R756 avss.t275 avss.n112 59.46
R757 avss.t110 avss.n109 59.46
R758 avss.t217 avss.n106 59.46
R759 avss.t132 avss.n103 59.46
R760 avss.t159 avss.n100 59.46
R761 avss.t323 avss.n97 59.46
R762 avss.t290 avss.n94 59.46
R763 avss.t363 avss.n91 59.46
R764 avss.t180 avss.n88 59.46
R765 avss.t153 avss.n85 59.46
R766 avss.t329 avss.n82 59.46
R767 avss.t332 avss.n79 59.46
R768 avss.t137 avss.n76 59.46
R769 avss.t189 avss.n73 59.46
R770 avss.t277 avss.n70 59.46
R771 avss.t84 avss.t157 59.3854
R772 avss.t365 avss.t102 58.5371
R773 avss.t188 avss.t130 57.6887
R774 avss.n644 avss.t13 57.0602
R775 avss.n763 avss.t172 56.675
R776 avss.t103 avss.t12 55.1437
R777 avss.t298 avss.t186 54.4857
R778 avss.t272 avss.t322 54.2953
R779 avss.t341 avss.t306 53.4469
R780 avss.n589 avss.n554 53.1823
R781 avss.n589 avss.n562 53.1823
R782 avss.n617 avss.n552 53.1823
R783 avss.n618 avss.n617 53.1823
R784 avss.n373 avss.n371 53.1823
R785 avss.n763 avss.n371 53.1823
R786 avss.n770 avss.n372 53.1823
R787 avss.n763 avss.n372 53.1823
R788 avss.n18 avss.t158 52.9509
R789 avss.t259 avss.n8 52.5315
R790 avss.n46 avss.t89 51.9277
R791 avss.t113 avss.t249 50.0535
R792 avss.n623 avss.n622 49.8123
R793 avss.n586 avss.n585 49.8123
R794 avss.n757 avss.n755 49.8123
R795 avss.n759 avss.n381 49.8123
R796 avss.t30 avss.t119 49.2052
R797 avss.t42 avss.n409 48.6621
R798 avss.t135 avss.t156 48.3568
R799 avss.n673 avss.t267 47.2902
R800 avss.t128 avss.t334 45.8117
R801 avss.t292 avss.t319 45.5327
R802 avss.t54 avss.t320 45.5327
R803 avss.t10 avss.t198 45.5327
R804 avss.n11 avss.n9 45.0005
R805 avss.t89 avss.n9 45.0005
R806 avss.n876 avss.n10 45.0005
R807 avss.t89 avss.n10 45.0005
R808 avss.t129 avss.t52 44.9634
R809 avss.n764 avss.t235 44.1554
R810 avss.n762 avss.t174 44.1554
R811 avss.t215 avss.t274 44.115
R812 avss.t326 avss.n18 43.7421
R813 avss.n343 avss.t109 43.6909
R814 avss.t136 avss.n342 43.6909
R815 avss.n419 avss.n410 43.3803
R816 avss.n428 avss.n404 43.3803
R817 avss.n422 avss.n410 43.3803
R818 avss.n428 avss.n427 43.3803
R819 avss.t114 avss.n49 42.7523
R820 avss.n859 avss.n858 42.7189
R821 avss.n774 avss.n370 42.3223
R822 avss.t199 avss.t298 42.2073
R823 avss.t273 avss.t214 40.7216
R824 avss.t288 avss.t250 39.8732
R825 avss.n774 avss.t174 39.7462
R826 avss.t65 avss.t257 39.0249
R827 avss.n794 avss.n793 38.6099
R828 avss.n794 avss.n53 38.6076
R829 avss.n793 avss.n792 38.5956
R830 avss.t257 avss.t136 36.4798
R831 avss.t314 avss.n879 36.324
R832 avss.n318 avss.n311 36.1417
R833 avss.n312 avss.n311 36.1417
R834 avss.n299 avss.n72 36.1417
R835 avss.n305 avss.n72 36.1417
R836 avss.n287 avss.n75 36.1417
R837 avss.n294 avss.n75 36.1417
R838 avss.n275 avss.n78 36.1417
R839 avss.n282 avss.n78 36.1417
R840 avss.n263 avss.n81 36.1417
R841 avss.n270 avss.n81 36.1417
R842 avss.n251 avss.n84 36.1417
R843 avss.n258 avss.n84 36.1417
R844 avss.n239 avss.n87 36.1417
R845 avss.n246 avss.n87 36.1417
R846 avss.n227 avss.n90 36.1417
R847 avss.n234 avss.n90 36.1417
R848 avss.n215 avss.n93 36.1417
R849 avss.n222 avss.n93 36.1417
R850 avss.n203 avss.n96 36.1417
R851 avss.n210 avss.n96 36.1417
R852 avss.n191 avss.n99 36.1417
R853 avss.n198 avss.n99 36.1417
R854 avss.n179 avss.n102 36.1417
R855 avss.n186 avss.n102 36.1417
R856 avss.n167 avss.n105 36.1417
R857 avss.n174 avss.n105 36.1417
R858 avss.n155 avss.n108 36.1417
R859 avss.n162 avss.n108 36.1417
R860 avss.n143 avss.n111 36.1417
R861 avss.n150 avss.n111 36.1417
R862 avss.n131 avss.n114 36.1417
R863 avss.n138 avss.n114 36.1417
R864 avss.n120 avss.n119 36.1417
R865 avss.n126 avss.n120 36.1417
R866 avss.n338 avss.n62 36.1417
R867 avss.n791 avss.n53 35.7393
R868 avss.t250 avss.t289 35.6315
R869 avss.n420 avss.n418 35.5561
R870 avss.n415 avss.n412 35.5561
R871 avss.n487 avss.n476 35.1094
R872 avss.n533 avss.n454 35.1094
R873 avss.t214 avss.t78 34.7831
R874 avss.n340 avss.n339 34.4123
R875 avss.n341 avss.n340 34.4123
R876 avss.n345 avss.n344 34.4123
R877 avss.n344 avss.n343 34.4123
R878 avss.n801 avss.t304 33.2544
R879 avss.n650 avss.n22 32.5005
R880 avss.t115 avss.n650 32.5005
R881 avss.n648 avss.n636 32.5005
R882 avss.n636 avss.t14 32.5005
R883 avss.n649 avss.n637 32.5005
R884 avss.n637 avss.t14 32.5005
R885 avss.n878 avss.n877 32.5005
R886 avss.n879 avss.n878 32.5005
R887 avss.n875 avss.n874 32.5005
R888 avss.n874 avss.n873 32.5005
R889 avss.n871 avss.n870 32.5005
R890 avss.n872 avss.n871 32.5005
R891 avss.n861 avss.n860 32.5005
R892 avss.n860 avss.n859 32.5005
R893 avss.n857 avss.n856 32.5005
R894 avss.n858 avss.n857 32.5005
R895 avss.n342 avss.t135 31.8139
R896 avss.n859 avss.t151 31.4638
R897 avss.t20 avss.t215 31.3897
R898 avss.t325 avss.t129 30.5413
R899 avss.t331 avss.t128 29.693
R900 avss.n494 avss.n471 29.6559
R901 avss.n511 avss.n510 29.6559
R902 avss.n527 avss.n526 29.6559
R903 avss.n416 avss.n407 29.4328
R904 avss.n413 avss.n408 29.4328
R905 avss.n414 avss.n407 29.4328
R906 avss.n408 avss.n405 29.4328
R907 avss.n677 avss.n676 28.9887
R908 avss.n768 avss.n366 28.9887
R909 avss.t99 avss.t54 28.9058
R910 avss.t82 avss.t143 28.65
R911 avss.t156 avss.t28 27.1479
R912 avss.n649 avss.n639 27.1064
R913 avss.n648 avss.n638 27.1064
R914 avss.n538 avss.n537 26.8634
R915 avss.t108 avss.t16 26.5545
R916 avss.n819 avss.t57 26.4633
R917 avss.n814 avss.t33 26.4633
R918 avss.n41 avss.t48 26.4633
R919 avss.n809 avss.t66 26.4633
R920 avss.n828 avss.t93 26.4633
R921 avss.n834 avss.t4 26.4633
R922 avss.n844 avss.t90 26.4633
R923 avss.n839 avss.t96 26.4633
R924 avss.n28 avss.t15 26.4633
R925 avss.n36 avss.t37 26.4633
R926 avss.t119 avss.t362 26.2995
R927 avss.t201 avss.t317 26.092
R928 avss.t249 avss.t112 25.4512
R929 avss.n645 avss.t35 25.2191
R930 avss.n642 avss.t68 25.2191
R931 avss.t89 avss.t199 23.7898
R932 avss.n16 avss.t316 23.7186
R933 avss.n864 avss.t197 23.4728
R934 avss.n867 avss.t318 23.4728
R935 avss.n16 avss.t299 23.4728
R936 avss.t185 avss.t82 23.2782
R937 avss.n858 avss.t304 22.5108
R938 avss.n676 avss.n675 22.5005
R939 avss.n675 avss.n674 22.5005
R940 avss.n561 avss.n560 22.5005
R941 avss.n674 avss.n561 22.5005
R942 avss.n366 avss.n364 22.5005
R943 avss.n377 avss.n364 22.5005
R944 avss.n777 avss.n365 22.5005
R945 avss.n377 avss.n365 22.5005
R946 avss.n872 avss.t252 22.255
R947 avss.t320 avss.t185 22.255
R948 avss.n765 avss.t247 22.0815
R949 avss.t305 avss.t341 22.0578
R950 avss.n629 avss.n567 21.3347
R951 avss.t76 avss.t272 21.2094
R952 avss.n629 avss.n628 21.1018
R953 avss.n628 avss.n627 20.9741
R954 avss.n622 avss.n621 20.8934
R955 avss.n621 avss.n620 20.8934
R956 avss.n587 avss.n586 20.8934
R957 avss.n588 avss.n587 20.8934
R958 avss.n757 avss.n756 20.8934
R959 avss.n756 avss.n376 20.8934
R960 avss.n760 avss.n759 20.8934
R961 avss.n761 avss.n760 20.8934
R962 avss.t196 avss.t141 20.7202
R963 avss.n818 avss.n817 20.3733
R964 avss.n816 avss.n815 20.3733
R965 avss.n806 avss.n805 20.3733
R966 avss.n808 avss.n807 20.3733
R967 avss.n831 avss.n830 20.3733
R968 avss.n833 avss.n832 20.3733
R969 avss.n843 avss.n842 20.3733
R970 avss.n841 avss.n840 20.3733
R971 avss.n33 avss.n32 20.3733
R972 avss.n35 avss.n34 20.3733
R973 avss.t327 avss.t103 20.361
R974 avss avss.n424 20.2672
R975 avss.n14 avss.n12 20.1729
R976 avss.n18 avss.n12 20.1729
R977 avss.n15 avss.n13 20.1729
R978 avss.n18 avss.n13 20.1729
R979 avss.n866 avss.n865 20.1668
R980 avss.t239 avss.n764 19.7448
R981 avss.t172 avss.n762 19.7448
R982 avss.n349 avss.t313 19.4214
R983 avss.t258 avss.n341 18.2402
R984 avss.n819 avss.t59 18.0193
R985 avss.t34 avss.n814 18.0193
R986 avss.n41 avss.t50 18.0193
R987 avss.n809 avss.t67 18.0193
R988 avss.n828 avss.t95 18.0193
R989 avss.n834 avss.t6 18.0193
R990 avss.n844 avss.t92 18.0193
R991 avss.t97 avss.n839 18.0193
R992 avss.n28 avss.t18 18.0193
R993 avss.n36 avss.t38 18.0193
R994 avss.n517 avss.n516 17.9618
R995 avss.n504 avss.n468 17.9618
R996 avss.n504 avss.n503 17.9618
R997 avss.n516 avss.n464 17.9618
R998 avss.n431 avss.n430 17.9561
R999 avss.t130 avss.t187 17.816
R1000 avss.n626 avss.n566 17.6946
R1001 avss.n431 avss.n402 17.6005
R1002 avss.n645 avss.t36 17.2863
R1003 avss.n642 avss.t69 17.2863
R1004 avss.t102 avss.t8 16.9676
R1005 avss.n484 avss 16.7292
R1006 avss.t319 avss.t99 16.6274
R1007 avss.n572 avss.t353 16.5305
R1008 avss.n572 avss.t345 16.5305
R1009 avss.n570 avss.t347 16.5305
R1010 avss.n570 avss.t351 16.5305
R1011 avss.n576 avss.t349 16.5305
R1012 avss.n576 avss.t355 16.5305
R1013 avss.n574 avss.t343 16.5305
R1014 avss.n574 avss.t359 16.5305
R1015 avss.n545 avss.t232 16.5305
R1016 avss.n545 avss.t71 16.5305
R1017 avss.n543 avss.t285 16.5305
R1018 avss.n543 avss.t62 16.5305
R1019 avss.n549 avss.t228 16.5305
R1020 avss.n549 avss.t226 16.5305
R1021 avss.n611 avss.t283 16.5305
R1022 avss.n611 avss.t286 16.5305
R1023 avss.t47 avss.n595 16.5305
R1024 avss.n595 avss.t230 16.5305
R1025 avss.n608 avss.t41 16.5305
R1026 avss.n608 avss.t284 16.5305
R1027 avss.n385 avss.t244 16.5305
R1028 avss.n385 avss.t238 16.5305
R1029 avss.n383 avss.t234 16.5305
R1030 avss.n383 avss.t246 16.5305
R1031 avss.n389 avss.t248 16.5305
R1032 avss.n389 avss.t240 16.5305
R1033 avss.n387 avss.t236 16.5305
R1034 avss.n387 avss.t173 16.5305
R1035 avss.n711 avss.t338 16.5305
R1036 avss.n711 avss.t86 16.5305
R1037 avss.n709 avss.t126 16.5305
R1038 avss.n709 avss.t25 16.5305
R1039 avss.n395 avss.t337 16.5305
R1040 avss.n395 avss.t340 16.5305
R1041 avss.n393 avss.t125 16.5305
R1042 avss.n393 avss.t124 16.5305
R1043 avss.n748 avss.t3 16.5305
R1044 avss.n748 avss.t339 16.5305
R1045 avss.n745 avss.t45 16.5305
R1046 avss.n745 avss.t127 16.5305
R1047 avss.t157 avss.t216 16.1193
R1048 avss.n627 avss.n625 15.8429
R1049 avss.n425 avss 15.2894
R1050 avss.n855 avss.n17 14.9605
R1051 avss.n869 avss.n868 14.9605
R1052 avss.n863 avss.n862 14.9605
R1053 avss.n853 avss.n852 14.9605
R1054 avss.t163 avss.t326 14.8368
R1055 avss.t141 avss.t179 14.581
R1056 avss.n688 avss.t70 14.0925
R1057 avss.n540 avss.t60 14.0925
R1058 avss.n596 avss.t46 14.0925
R1059 avss.n607 avss.t39 14.0925
R1060 avss.n747 avss.t1 14.0925
R1061 avss.n744 avss.t44 14.0925
R1062 avss.n719 avss.t85 14.0925
R1063 avss.n706 avss.t23 14.0925
R1064 avss.n46 avss.t315 14.0694
R1065 avss.t143 avss.n798 13.0463
R1066 avss.n479 avss 12.9272
R1067 avss.n873 avss.t186 12.7905
R1068 avss.n21 avss.n19 12.7179
R1069 avss.t282 avss.n19 12.7179
R1070 avss.n854 avss.n20 12.7179
R1071 avss.t282 avss.n20 12.7179
R1072 avss.t170 avss.n376 12.513
R1073 avss.n880 avss.t212 12.2789
R1074 avss.n358 avss.n355 12.189
R1075 avss.n421 avss.n420 12.0894
R1076 avss.n418 avss.n417 12.0894
R1077 avss.n426 avss.n402 12.0894
R1078 avss.n430 avss.n403 12.0894
R1079 avss.n656 avss.t209 11.9874
R1080 avss.t161 avss.t176 11.8775
R1081 avss.n888 avss.n887 11.8447
R1082 avss.n362 avss.t16 11.7601
R1083 avss.n377 avss.t170 11.409
R1084 avss.t32 avss.t336 11.0291
R1085 avss.n368 avss.n49 10.9999
R1086 avss.n765 avss.n376 10.673
R1087 avss.n392 avss.n381 10.3632
R1088 avss.n755 avss.n754 10.3105
R1089 avss.n624 avss.n623 10.3105
R1090 avss.n585 avss.n584 10.3105
R1091 avss.n822 avss.n804 9.42076
R1092 avss.n812 avss.n804 9.42076
R1093 avss.n352 avss.n57 9.35869
R1094 avss.n351 avss.n58 9.35222
R1095 avss.n350 avss.n59 9.34791
R1096 avss.n353 avss.n56 9.33929
R1097 avss.n354 avss.n55 9.33929
R1098 avss.n317 avss.n316 9.30641
R1099 avss.n316 avss.n315 9.3005
R1100 avss.n318 avss.n317 9.3005
R1101 avss.n314 avss.n311 9.3005
R1102 avss.n313 avss.n312 9.3005
R1103 avss.n666 avss.n639 9.3005
R1104 avss.n640 avss.n638 9.3005
R1105 avss.n654 avss.n653 9.3005
R1106 avss.n786 avss.n357 9.3005
R1107 avss.n124 avss.n123 9.3005
R1108 avss.n123 avss.n122 9.3005
R1109 avss.n136 avss.n135 9.3005
R1110 avss.n135 avss.n134 9.3005
R1111 avss.n148 avss.n147 9.3005
R1112 avss.n147 avss.n146 9.3005
R1113 avss.n160 avss.n159 9.3005
R1114 avss.n159 avss.n158 9.3005
R1115 avss.n172 avss.n171 9.3005
R1116 avss.n171 avss.n170 9.3005
R1117 avss.n184 avss.n183 9.3005
R1118 avss.n183 avss.n182 9.3005
R1119 avss.n196 avss.n195 9.3005
R1120 avss.n195 avss.n194 9.3005
R1121 avss.n208 avss.n207 9.3005
R1122 avss.n207 avss.n206 9.3005
R1123 avss.n220 avss.n219 9.3005
R1124 avss.n219 avss.n218 9.3005
R1125 avss.n232 avss.n231 9.3005
R1126 avss.n231 avss.n230 9.3005
R1127 avss.n244 avss.n243 9.3005
R1128 avss.n243 avss.n242 9.3005
R1129 avss.n256 avss.n255 9.3005
R1130 avss.n255 avss.n254 9.3005
R1131 avss.n268 avss.n267 9.3005
R1132 avss.n267 avss.n266 9.3005
R1133 avss.n280 avss.n279 9.3005
R1134 avss.n279 avss.n278 9.3005
R1135 avss.n292 avss.n291 9.3005
R1136 avss.n291 avss.n290 9.3005
R1137 avss.n302 avss.n0 9.3005
R1138 avss.n303 avss.n302 9.3005
R1139 avss.n132 avss.n131 9.3005
R1140 avss.n133 avss.n114 9.3005
R1141 avss.n138 avss.n137 9.3005
R1142 avss.n144 avss.n143 9.3005
R1143 avss.n145 avss.n111 9.3005
R1144 avss.n150 avss.n149 9.3005
R1145 avss.n156 avss.n155 9.3005
R1146 avss.n157 avss.n108 9.3005
R1147 avss.n162 avss.n161 9.3005
R1148 avss.n168 avss.n167 9.3005
R1149 avss.n169 avss.n105 9.3005
R1150 avss.n174 avss.n173 9.3005
R1151 avss.n180 avss.n179 9.3005
R1152 avss.n181 avss.n102 9.3005
R1153 avss.n186 avss.n185 9.3005
R1154 avss.n192 avss.n191 9.3005
R1155 avss.n193 avss.n99 9.3005
R1156 avss.n198 avss.n197 9.3005
R1157 avss.n204 avss.n203 9.3005
R1158 avss.n205 avss.n96 9.3005
R1159 avss.n210 avss.n209 9.3005
R1160 avss.n216 avss.n215 9.3005
R1161 avss.n217 avss.n93 9.3005
R1162 avss.n222 avss.n221 9.3005
R1163 avss.n228 avss.n227 9.3005
R1164 avss.n229 avss.n90 9.3005
R1165 avss.n234 avss.n233 9.3005
R1166 avss.n240 avss.n239 9.3005
R1167 avss.n241 avss.n87 9.3005
R1168 avss.n246 avss.n245 9.3005
R1169 avss.n252 avss.n251 9.3005
R1170 avss.n253 avss.n84 9.3005
R1171 avss.n258 avss.n257 9.3005
R1172 avss.n264 avss.n263 9.3005
R1173 avss.n265 avss.n81 9.3005
R1174 avss.n270 avss.n269 9.3005
R1175 avss.n276 avss.n275 9.3005
R1176 avss.n277 avss.n78 9.3005
R1177 avss.n282 avss.n281 9.3005
R1178 avss.n288 avss.n287 9.3005
R1179 avss.n289 avss.n75 9.3005
R1180 avss.n294 avss.n293 9.3005
R1181 avss.n300 avss.n299 9.3005
R1182 avss.n301 avss.n72 9.3005
R1183 avss.n305 avss.n304 9.3005
R1184 avss.n119 avss.n60 9.3005
R1185 avss.n121 avss.n120 9.3005
R1186 avss.n126 avss.n125 9.3005
R1187 avss.n347 avss.n346 9.3005
R1188 avss.n789 avss.n788 9.20927
R1189 avss.t237 avss.n377 8.83289
R1190 avss.t235 avss.n763 8.83289
R1191 avss.n657 avss.n655 8.81442
R1192 avss.n604 avss.t393 8.80038
R1193 avss.n603 avss.t382 8.80038
R1194 avss.n602 avss.t375 8.80038
R1195 avss.n601 avss.t397 8.80038
R1196 avss.n600 avss.t377 8.80038
R1197 avss.n599 avss.t366 8.80038
R1198 avss.n598 avss.t387 8.80038
R1199 avss.n539 avss.t380 8.80038
R1200 avss.n741 avss.t376 8.80038
R1201 avss.n740 avss.t379 8.80038
R1202 avss.n739 avss.t386 8.80038
R1203 avss.n738 avss.t369 8.80038
R1204 avss.n737 avss.t384 8.80038
R1205 avss.n736 avss.t396 8.80038
R1206 avss.n735 avss.t374 8.80038
R1207 avss.n734 avss.t381 8.80038
R1208 avss.n694 avss.t383 8.73382
R1209 avss.n695 avss.t372 8.73382
R1210 avss.n696 avss.t367 8.73382
R1211 avss.n697 avss.t389 8.73382
R1212 avss.n698 avss.t368 8.73382
R1213 avss.n699 avss.t390 8.73382
R1214 avss.n700 avss.t373 8.73382
R1215 avss.n701 avss.t371 8.73382
R1216 avss.n725 avss.t388 8.73382
R1217 avss.n726 avss.t391 8.73382
R1218 avss.n727 avss.t395 8.73382
R1219 avss.n728 avss.t378 8.73382
R1220 avss.n729 avss.t394 8.73382
R1221 avss.n730 avss.t370 8.73382
R1222 avss.n731 avss.t385 8.73382
R1223 avss.n732 avss.t392 8.73382
R1224 avss.n492 avss.n475 8.61832
R1225 avss.n493 avss.n492 8.61832
R1226 avss.n494 avss.n493 8.61832
R1227 avss.n500 avss.n471 8.61832
R1228 avss.n501 avss.n500 8.61832
R1229 avss.n502 avss.n501 8.61832
R1230 avss.n509 avss.n467 8.61832
R1231 avss.n510 avss.n509 8.61832
R1232 avss.n511 avss.n465 8.61832
R1233 avss.n518 avss.n465 8.61832
R1234 avss.n460 avss.n452 8.61832
R1235 avss.n528 avss.n460 8.61832
R1236 avss.n528 avss.n527 8.61832
R1237 avss.n526 avss.n461 8.61832
R1238 avss.n520 avss.n461 8.61832
R1239 avss.n520 avss.n519 8.61832
R1240 avss.n486 avss.n485 8.61832
R1241 avss.n485 avss.n484 8.61832
R1242 avss.n479 avss.n451 8.61832
R1243 avss.t178 avss.t280 8.48406
R1244 avss.n655 avss.n358 8.4666
R1245 avss.n666 avss.n665 8.37766
R1246 avss.n665 avss.n640 8.37766
R1247 avss.n38 avss.n30 8.11041
R1248 avss.n848 avss.n30 8.11041
R1249 avss.n786 avss.n785 8.02619
R1250 avss.n785 avss.n358 8.00675
R1251 avss.n667 avss.n640 7.938
R1252 avss.n667 avss.n666 7.938
R1253 avss.t192 avss.t182 7.63571
R1254 avss.n702 avss.n539 7.62598
R1255 avss.n734 avss.n733 7.62598
R1256 avss.n658 avss.n654 7.48375
R1257 avss.n424 avss.n421 7.46717
R1258 avss.n426 avss.n425 7.46717
R1259 avss.n417 avss.n415 7.46717
R1260 avss.n412 avss.n403 7.46717
R1261 avss.n658 avss.n657 7.16066
R1262 avss.t315 avss.t204 6.90708
R1263 avss.n654 avss.n356 6.89147
R1264 avss.n786 avss.n356 6.89083
R1265 avss.n48 avss.n45 6.88285
R1266 avss.n362 avss.n48 6.88285
R1267 avss.n47 avss.n44 6.88285
R1268 avss.n47 avss.n46 6.88285
R1269 avss.t310 avss.t74 6.78735
R1270 avss.n669 avss.n668 6.5005
R1271 avss.n670 avss.n669 6.5005
R1272 avss.n664 avss.n663 6.5005
R1273 avss.n663 avss.n662 6.5005
R1274 avss.n680 avss.n551 6.47706
R1275 avss.n680 avss.n547 6.47706
R1276 avss.n613 avss.n610 6.47706
R1277 avss.n613 avss.n542 6.47706
R1278 avss.n750 avss.n375 6.47706
R1279 avss.n713 avss.n375 6.47706
R1280 avss.n401 avss.n374 6.47706
R1281 avss.n708 avss.n374 6.47706
R1282 avss.n535 avss.n451 6.46387
R1283 avss.n890 avss.n889 6.05765
R1284 avss.n800 avss.n799 5.90959
R1285 avss.n801 avss.n800 5.90959
R1286 avss.n803 avss.n802 5.90959
R1287 avss.n802 avss.n801 5.90959
R1288 avss.n368 avss.t10 5.88388
R1289 avss.n625 avss.n624 5.79451
R1290 avss.n889 avss.n2 5.78505
R1291 avss.n656 avss.n647 5.7846
R1292 avss.n646 avss.n645 5.76099
R1293 avss.n643 avss.n642 5.76099
R1294 avss.n813 avss.n812 5.70305
R1295 avss.n811 avss.n810 5.70305
R1296 avss.n836 avss.n835 5.70305
R1297 avss.n838 avss.n837 5.70305
R1298 avss.n38 avss.n37 5.70305
R1299 avss.n641 avss.n640 5.6605
R1300 avss.n820 avss.n819 5.6605
R1301 avss.n814 avss.n813 5.6605
R1302 avss.n822 avss.n821 5.6605
R1303 avss.n42 avss.n41 5.6605
R1304 avss.n810 avss.n809 5.6605
R1305 avss.n824 avss.n823 5.6605
R1306 avss.n829 avss.n828 5.6605
R1307 avss.n835 avss.n834 5.6605
R1308 avss.n827 avss.n31 5.6605
R1309 avss.n845 avss.n844 5.6605
R1310 avss.n839 avss.n838 5.6605
R1311 avss.n847 avss.n846 5.6605
R1312 avss.n29 avss.n28 5.6605
R1313 avss.n37 avss.n36 5.6605
R1314 avss.n849 avss.n848 5.6605
R1315 avss.n666 avss.n647 5.6605
R1316 avss.t158 avss.t165 5.62808
R1317 avss.n625 avss.n567 5.46789
R1318 avss.n630 avss.n565 5.27077
R1319 avss.n565 avss.n564 5.27077
R1320 avss.n566 avss.n563 5.27077
R1321 avss.n564 avss.n563 5.27077
R1322 avss.n784 avss.n783 5.27077
R1323 avss.n783 avss.n782 5.27077
R1324 avss.n660 avss.n659 5.27077
R1325 avss.n661 avss.n660 5.27077
R1326 avss.n544 avss.n542 5.07277
R1327 avss.n613 avss.n612 5.07277
R1328 avss.n610 avss.n609 5.07277
R1329 avss.n710 avss.n708 5.07277
R1330 avss.n394 avss.n374 5.07277
R1331 avss.n746 avss.n401 5.07277
R1332 avss.n632 avss.n631 5.0436
R1333 avss.n633 avss.n632 5.0436
R1334 avss.n569 avss.n568 5.0436
R1335 avss.n361 avss.n359 5.0436
R1336 avss.t108 avss.n361 5.0436
R1337 avss.n652 avss.n360 5.0436
R1338 avss.t108 avss.n360 5.0436
R1339 avss.n797 avss.n796 5.0436
R1340 avss.n798 avss.n797 5.0436
R1341 avss.n66 avss.n54 5.0436
R1342 avss.n67 avss.n66 5.0436
R1343 avss.n447 avss.n446 5.0005
R1344 avss.n446 avss.n445 5.0005
R1345 avss.n438 avss.n434 5.0005
R1346 avss.n444 avss.n438 5.0005
R1347 avss.n442 avss.n441 5.0005
R1348 avss.n443 avss.n442 5.0005
R1349 avss.n440 avss.n437 5.0005
R1350 avss.n439 avss.n437 5.0005
R1351 avss.n547 avss.n546 4.95167
R1352 avss.n592 avss.n551 4.95167
R1353 avss.n713 avss.n712 4.95167
R1354 avss.n750 avss.n749 4.95167
R1355 avss.n791 avss.n790 4.86769
R1356 avss.n63 avss.n62 4.6805
R1357 avss.t30 avss.n63 4.6805
R1358 avss.n65 avss.n64 4.6805
R1359 avss.t30 avss.n65 4.6805
R1360 avss.n733 avss.n732 4.60905
R1361 avss.n702 avss.n701 4.60905
R1362 avss.n541 avss.n540 4.5005
R1363 avss.n689 avss.n688 4.5005
R1364 avss.n681 avss.n680 4.5005
R1365 avss.n691 avss.n690 4.5005
R1366 avss.n693 avss.n692 4.5005
R1367 avss.n607 avss.n606 4.5005
R1368 avss.n597 avss.n596 4.5005
R1369 avss.n605 avss.n591 4.5005
R1370 avss.n594 avss.n593 4.5005
R1371 avss.n397 avss.n375 4.5005
R1372 avss.n707 avss.n706 4.5005
R1373 avss.n720 avss.n719 4.5005
R1374 avss.n724 avss.n723 4.5005
R1375 avss.n722 avss.n721 4.5005
R1376 avss.n744 avss.n743 4.5005
R1377 avss.n747 avss.n399 4.5005
R1378 avss.n742 avss.n400 4.5005
R1379 avss.n752 avss.n751 4.5005
R1380 avss.n435 avss.n432 4.3603
R1381 avss.n449 avss.n433 4.34678
R1382 avss.n435 avss.n433 4.34003
R1383 avss.n641 avss.n26 4.00655
R1384 avss.n616 avss.n614 3.9532
R1385 avss.n616 avss.n615 3.9532
R1386 avss.n679 avss.n553 3.9532
R1387 avss.n615 avss.n553 3.9532
R1388 avss.n767 avss.n766 3.9532
R1389 avss.n766 avss.n765 3.9532
R1390 avss.n773 avss.n772 3.9532
R1391 avss.n774 avss.n773 3.9532
R1392 avss.n889 avss.n888 3.94537
R1393 avss.n704 avss.n703 3.9105
R1394 avss.n798 avss.t198 3.83749
R1395 avss.n450 avss.n449 3.78259
R1396 avss.n594 avss.n548 3.77378
R1397 avss.n753 avss.n752 3.77378
R1398 avss.n682 avss.n681 3.77209
R1399 avss.n398 avss.n397 3.77209
R1400 avss.n690 avss.n687 3.77014
R1401 avss.n721 avss.n718 3.77014
R1402 avss.n852 avss.n851 3.68964
R1403 avss.n821 avss.n40 3.57087
R1404 avss.n825 avss.n824 3.57087
R1405 avss.n827 avss.n826 3.57087
R1406 avss.n846 avss.n27 3.57087
R1407 avss.n850 avss.n849 3.57087
R1408 avss.n392 avss.n391 3.4105
R1409 avss.n717 avss.n716 3.4105
R1410 avss.n686 avss.n685 3.4105
R1411 avss.n579 avss.n578 3.4105
R1412 avss.n817 avss.t147 3.3065
R1413 avss.n817 avss.t58 3.3065
R1414 avss.n815 avss.t34 3.3065
R1415 avss.n815 avss.t146 3.3065
R1416 avss.n805 avss.t261 3.3065
R1417 avss.n805 avss.t49 3.3065
R1418 avss.t67 avss.n808 3.3065
R1419 avss.n808 avss.t148 3.3065
R1420 avss.n830 avss.t144 3.3065
R1421 avss.n830 avss.t94 3.3065
R1422 avss.t6 avss.n833 3.3065
R1423 avss.n833 avss.t142 3.3065
R1424 avss.n842 avss.t149 3.3065
R1425 avss.n842 avss.t91 3.3065
R1426 avss.n840 avss.t97 3.3065
R1427 avss.n840 avss.t262 3.3065
R1428 avss.n32 avss.t145 3.3065
R1429 avss.n32 avss.t17 3.3065
R1430 avss.t38 avss.n35 3.3065
R1431 avss.n35 avss.t260 3.3065
R1432 avss.n865 avss.t166 3.3065
R1433 avss.n865 avss.t164 3.3065
R1434 avss.t115 avss.n651 3.2875
R1435 avss.n593 avss.n551 3.23878
R1436 avss.n691 avss.n547 3.23878
R1437 avss.n610 avss.n591 3.23878
R1438 avss.n692 avss.n542 3.23878
R1439 avss.n751 avss.n750 3.23878
R1440 avss.n722 avss.n713 3.23878
R1441 avss.n401 avss.n400 3.23878
R1442 avss.n723 avss.n708 3.23878
R1443 avss.n733 avss.n705 3.22196
R1444 avss.n694 avss.n693 3.21858
R1445 avss.n725 avss.n724 3.21858
R1446 avss.n605 avss.n604 3.12292
R1447 avss.n742 avss.n741 3.12292
R1448 avss.n536 avss.n535 3.1005
R1449 avss.n68 avss.t255 2.96975
R1450 avss.n792 avss.n791 2.83532
R1451 avss.n887 avss.n3 2.6005
R1452 avss.t131 avss.t0 2.54557
R1453 avss.n848 avss.n847 2.42291
R1454 avss.n847 avss.n31 2.42291
R1455 avss.n823 avss.n822 2.42291
R1456 avss.n812 avss.n811 2.42291
R1457 avss.n837 avss.n836 2.42291
R1458 avss.n837 avss.n38 2.42291
R1459 avss.n502 avss.n467 2.40842
R1460 avss.n519 avss.n518 2.40842
R1461 avss.n537 avss.n431 2.32925
R1462 avss.n787 avss.n786 2.31886
R1463 avss.n654 avss.n26 2.31886
R1464 avss.n486 avss.n475 2.28169
R1465 avss.n534 avss.n452 2.28169
R1466 avss.n705 avss.n704 2.28019
R1467 avss.n440 avss.n436 2.25932
R1468 avss.n657 avss.n656 2.2505
R1469 avss.n704 avss.n355 2.221
R1470 avss.n536 avss.n450 2.17339
R1471 avss.n535 avss.n534 2.15496
R1472 avss.n703 avss.n702 2.12151
R1473 avss.n593 avss.n591 2.11769
R1474 avss.n692 avss.n691 2.11769
R1475 avss.n751 avss.n400 2.11769
R1476 avss.n723 avss.n722 2.11769
R1477 avss.n788 avss.n355 2.058
R1478 avss.n703 avss.n538 1.90581
R1479 avss.n686 avss.n538 1.80585
R1480 avss.n823 avss.n43 1.80222
R1481 avss.n811 avss.n39 1.80222
R1482 avss.t152 avss.t208 1.69721
R1483 avss.n352 avss.n351 1.6605
R1484 avss.n753 avss.n398 1.58008
R1485 avss.n718 avss.n398 1.58008
R1486 avss.n687 avss.n682 1.58008
R1487 avss.n682 avss.n548 1.58008
R1488 avss.n795 avss.n51 1.50436
R1489 avss.n342 avss.n51 1.50436
R1490 avss.n52 avss.n50 1.50436
R1491 avss.n342 avss.n50 1.50436
R1492 avss.n348 avss.n60 1.48467
R1493 avss.n330 avss.n1 1.34141
R1494 avss.n351 avss.n350 1.338
R1495 avss.n347 avss.n61 1.32209
R1496 avss.n801 avss.t292 1.2795
R1497 avss.n354 avss.n353 1.27675
R1498 avss.t213 avss.n322 1.27303
R1499 avss.n651 avss.n363 1.27293
R1500 avss.n325 avss.n324 1.14936
R1501 avss.n335 avss.n334 1.14936
R1502 avss.n336 avss.n335 1.14839
R1503 avss.n324 avss.n323 1.14811
R1504 avss.n323 avss.n61 1.08686
R1505 avss.n326 avss.n325 1.08686
R1506 avss.n327 avss.n326 1.08686
R1507 avss.n329 avss.n328 1.08686
R1508 avss.n334 avss.n333 1.08686
R1509 avss.n333 avss.n332 1.08686
R1510 avss.n332 avss.n331 1.08686
R1511 avss.n331 avss.n330 1.08686
R1512 avss.n328 avss.n327 1.08005
R1513 avss.n818 avss.n816 1.05355
R1514 avss.n807 avss.n806 1.05355
R1515 avss.n832 avss.n831 1.05355
R1516 avss.n843 avss.n841 1.05355
R1517 avss.n34 avss.n33 1.05355
R1518 avss.n353 avss.n352 1.00987
R1519 avss.n337 avss.n336 1.00505
R1520 avss.n717 avss.n705 1.00226
R1521 avss.n646 avss.n644 0.955426
R1522 avss.n644 avss.n643 0.953203
R1523 avss.n789 avss.n1 0.902375
R1524 avss.n349 avss.n348 0.839875
R1525 avss.n604 avss.n603 0.807835
R1526 avss.n603 avss.n602 0.807835
R1527 avss.n602 avss.n601 0.807835
R1528 avss.n601 avss.n600 0.807835
R1529 avss.n600 avss.n599 0.807835
R1530 avss.n599 avss.n598 0.807835
R1531 avss.n598 avss.n539 0.807835
R1532 avss.n741 avss.n740 0.807835
R1533 avss.n740 avss.n739 0.807835
R1534 avss.n739 avss.n738 0.807835
R1535 avss.n738 avss.n737 0.807835
R1536 avss.n737 avss.n736 0.807835
R1537 avss.n736 avss.n735 0.807835
R1538 avss.n735 avss.n734 0.807835
R1539 avss.n695 avss.n694 0.80776
R1540 avss.n696 avss.n695 0.80776
R1541 avss.n697 avss.n696 0.80776
R1542 avss.n698 avss.n697 0.80776
R1543 avss.n699 avss.n698 0.80776
R1544 avss.n700 avss.n699 0.80776
R1545 avss.n701 avss.n700 0.80776
R1546 avss.n726 avss.n725 0.80776
R1547 avss.n727 avss.n726 0.80776
R1548 avss.n728 avss.n727 0.80776
R1549 avss.n729 avss.n728 0.80776
R1550 avss.n730 avss.n729 0.80776
R1551 avss.n731 avss.n730 0.80776
R1552 avss.n732 avss.n731 0.80776
R1553 avss.n891 avss.n890 0.79175
R1554 avss.n448 avss.n434 0.753441
R1555 avss.n577 avss.n575 0.695812
R1556 avss.n689 avss.n541 0.695812
R1557 avss.n546 avss.n544 0.695812
R1558 avss.n609 avss.n592 0.695812
R1559 avss.n606 avss.n597 0.695812
R1560 avss.n715 avss.n714 0.695812
R1561 avss.n390 avss.n388 0.695812
R1562 avss.n712 avss.n710 0.695812
R1563 avss.n396 avss.n394 0.695812
R1564 avss.n749 avss.n746 0.695812
R1565 avss.n720 avss.n707 0.695812
R1566 avss.n743 avss.n399 0.695812
R1567 avss.n684 avss.n683 0.695812
R1568 avss.t243 avss.n378 0.69443
R1569 avss.n573 avss.n571 0.679185
R1570 avss.n386 avss.n384 0.679185
R1571 avss.n612 avss.n550 0.676856
R1572 avss.n578 avss.n577 0.654797
R1573 avss.n391 avss.n390 0.654797
R1574 avss.n852 avss.n25 0.635318
R1575 avss.n43 avss.n31 0.62119
R1576 avss.n836 avss.n39 0.62119
R1577 avss.n693 avss.n541 0.572766
R1578 avss.n606 avss.n605 0.572766
R1579 avss.n724 avss.n707 0.572766
R1580 avss.n743 avss.n742 0.572766
R1581 avss.n450 avss.n432 0.571446
R1582 avss.n816 avss.n813 0.527027
R1583 avss.n820 avss.n818 0.527027
R1584 avss.n810 avss.n807 0.527027
R1585 avss.n806 avss.n42 0.527027
R1586 avss.n835 avss.n832 0.527027
R1587 avss.n831 avss.n829 0.527027
R1588 avss.n841 avss.n838 0.527027
R1589 avss.n845 avss.n843 0.527027
R1590 avss.n37 avss.n34 0.527027
R1591 avss.n33 avss.n29 0.527027
R1592 avss.t5 avss.n872 0.512098
R1593 avss.n851 avss.n26 0.505881
R1594 avss.n851 avss.n850 0.497189
R1595 avss.n850 avss.n27 0.478977
R1596 avss.n826 avss.n27 0.478977
R1597 avss.n826 avss.n825 0.478977
R1598 avss.n825 avss.n40 0.478977
R1599 avss.n690 avss.n689 0.451672
R1600 avss.n681 avss.n550 0.451672
R1601 avss.n597 avss.n594 0.451672
R1602 avss.n397 avss.n396 0.451672
R1603 avss.n721 avss.n720 0.451672
R1604 avss.n752 avss.n399 0.451672
R1605 avss.n788 avss.n787 0.387296
R1606 avss.n787 avss.n40 0.380881
R1607 avss.n890 avss.n1 0.364875
R1608 avss.n764 avss.t2 0.344476
R1609 avss.n716 avss.n715 0.311047
R1610 avss.n685 avss.n684 0.311047
R1611 avss.n867 avss.n866 0.291392
R1612 avss.n866 avss.n864 0.291392
R1613 avss.n436 avss.n435 0.274029
R1614 avss.n447 avss.n433 0.266214
R1615 avss.n449 avss.n448 0.266214
R1616 avss.n441 avss.n432 0.266214
R1617 avss.n132 avss 0.248811
R1618 avss.n144 avss 0.248811
R1619 avss.n156 avss 0.248811
R1620 avss.n168 avss 0.248811
R1621 avss.n180 avss 0.248811
R1622 avss.n192 avss 0.248811
R1623 avss.n204 avss 0.248811
R1624 avss.n216 avss 0.248811
R1625 avss.n228 avss 0.248811
R1626 avss.n240 avss 0.248811
R1627 avss.n252 avss 0.248811
R1628 avss.n264 avss 0.248811
R1629 avss.n276 avss 0.248811
R1630 avss.n288 avss 0.248811
R1631 avss.n300 avss 0.248811
R1632 avss.n718 avss.n717 0.237405
R1633 avss.n687 avss.n686 0.237405
R1634 avss.n23 avss.n17 0.182466
R1635 avss.n762 avss.t24 0.176117
R1636 avss.n350 avss.n349 0.153
R1637 avss.n348 avss.n347 0.128909
R1638 avss.n868 avss.n16 0.119588
R1639 avss.n754 avss.n753 0.118318
R1640 avss.n584 avss.n548 0.118318
R1641 avss.n45 avss.n43 0.11675
R1642 avss.n44 avss.n39 0.11675
R1643 avss.n24 avss.n23 0.11673
R1644 avss.n754 avss.n392 0.114189
R1645 avss.n584 avss.n579 0.114189
R1646 avss.n25 avss.n24 0.113554
R1647 avss.n668 avss.n667 0.109912
R1648 avss.n665 avss.n664 0.109912
R1649 avss avss.n891 0.107764
R1650 avss.n790 avss.n789 0.10175
R1651 avss.n799 avss.n30 0.0994362
R1652 avss.n804 avss.n803 0.0994362
R1653 avss.n627 avss.n626 0.0907913
R1654 avss.n659 avss.n658 0.0890714
R1655 avss.n785 avss.n784 0.0890714
R1656 avss.n630 avss.n629 0.0890714
R1657 avss.n652 avss.n356 0.0866111
R1658 avss.n793 avss.n54 0.0850455
R1659 avss.n796 avss.n53 0.0850455
R1660 avss.n655 avss.n359 0.0850455
R1661 avss.n628 avss.n569 0.0850455
R1662 avss.n631 avss.n567 0.0850455
R1663 avss.n337 avss.n329 0.0823182
R1664 avss.n314 avss.n313 0.0815811
R1665 avss.n121 avss.n60 0.0815811
R1666 avss.n133 avss.n132 0.0815811
R1667 avss.n145 avss.n144 0.0815811
R1668 avss.n157 avss.n156 0.0815811
R1669 avss.n169 avss.n168 0.0815811
R1670 avss.n181 avss.n180 0.0815811
R1671 avss.n193 avss.n192 0.0815811
R1672 avss.n205 avss.n204 0.0815811
R1673 avss.n217 avss.n216 0.0815811
R1674 avss.n229 avss.n228 0.0815811
R1675 avss.n241 avss.n240 0.0815811
R1676 avss.n253 avss.n252 0.0815811
R1677 avss.n265 avss.n264 0.0815811
R1678 avss.n277 avss.n276 0.0815811
R1679 avss.n289 avss.n288 0.0815811
R1680 avss.n301 avss.n300 0.0815811
R1681 avss.n338 avss.n337 0.0793136
R1682 avss.n537 avss.n536 0.0784703
R1683 avss.n680 avss.n679 0.0674065
R1684 avss.n614 avss.n613 0.0674065
R1685 avss.n772 avss.n374 0.0674065
R1686 avss.n767 avss.n375 0.0674065
R1687 avss.n125 avss.n122 0.0553986
R1688 avss.n137 avss.n134 0.0553986
R1689 avss.n149 avss.n146 0.0553986
R1690 avss.n161 avss.n158 0.0553986
R1691 avss.n173 avss.n170 0.0553986
R1692 avss.n185 avss.n182 0.0553986
R1693 avss.n197 avss.n194 0.0553986
R1694 avss.n209 avss.n206 0.0553986
R1695 avss.n221 avss.n218 0.0553986
R1696 avss.n233 avss.n230 0.0553986
R1697 avss.n245 avss.n242 0.0553986
R1698 avss.n257 avss.n254 0.0553986
R1699 avss.n269 avss.n266 0.0553986
R1700 avss.n281 avss.n278 0.0553986
R1701 avss.n293 avss.n290 0.0553986
R1702 avss.n304 avss.n303 0.0553986
R1703 avss.n863 avss.n17 0.0538514
R1704 avss.n624 avss.n579 0.0532162
R1705 avss.n891 avss 0.04675
R1706 avss.n647 avss.n646 0.0436892
R1707 avss.n821 avss.n820 0.0430541
R1708 avss.n824 avss.n42 0.0430541
R1709 avss.n829 avss.n827 0.0430541
R1710 avss.n846 avss.n845 0.0430541
R1711 avss.n849 avss.n29 0.0430541
R1712 avss.n868 avss.n867 0.0430541
R1713 avss.n643 avss.n641 0.0430541
R1714 avss.n864 avss.n863 0.0427365
R1715 avss.n313 avss 0.0410405
R1716 avss.n124 avss 0.0351284
R1717 avss.n136 avss 0.0351284
R1718 avss.n148 avss 0.0351284
R1719 avss.n160 avss 0.0351284
R1720 avss.n172 avss 0.0351284
R1721 avss.n184 avss 0.0351284
R1722 avss.n196 avss 0.0351284
R1723 avss.n208 avss 0.0351284
R1724 avss.n220 avss 0.0351284
R1725 avss.n232 avss 0.0351284
R1726 avss.n244 avss 0.0351284
R1727 avss.n256 avss 0.0351284
R1728 avss.n268 avss 0.0351284
R1729 avss.n280 avss 0.0351284
R1730 avss.n292 avss 0.0351284
R1731 avss avss.n0 0.0351284
R1732 avss.n315 avss.n2 0.0334392
R1733 avss.n315 avss.n314 0.0266824
R1734 avss.n122 avss.n121 0.0266824
R1735 avss.n134 avss.n133 0.0266824
R1736 avss.n146 avss.n145 0.0266824
R1737 avss.n158 avss.n157 0.0266824
R1738 avss.n170 avss.n169 0.0266824
R1739 avss.n182 avss.n181 0.0266824
R1740 avss.n194 avss.n193 0.0266824
R1741 avss.n206 avss.n205 0.0266824
R1742 avss.n218 avss.n217 0.0266824
R1743 avss.n230 avss.n229 0.0266824
R1744 avss.n242 avss.n241 0.0266824
R1745 avss.n254 avss.n253 0.0266824
R1746 avss.n266 avss.n265 0.0266824
R1747 avss.n278 avss.n277 0.0266824
R1748 avss.n290 avss.n289 0.0266824
R1749 avss.n303 avss.n301 0.0266824
R1750 avss.n792 avss.n52 0.0258406
R1751 avss.n795 avss.n794 0.0258406
R1752 avss.n317 avss.n2 0.0224595
R1753 avss.n578 avss.n573 0.0190811
R1754 avss.n391 avss.n386 0.0190811
R1755 avss.n125 avss.n124 0.00641216
R1756 avss.n137 avss.n136 0.00641216
R1757 avss.n149 avss.n148 0.00641216
R1758 avss.n161 avss.n160 0.00641216
R1759 avss.n173 avss.n172 0.00641216
R1760 avss.n185 avss.n184 0.00641216
R1761 avss.n197 avss.n196 0.00641216
R1762 avss.n209 avss.n208 0.00641216
R1763 avss.n221 avss.n220 0.00641216
R1764 avss.n233 avss.n232 0.00641216
R1765 avss.n245 avss.n244 0.00641216
R1766 avss.n257 avss.n256 0.00641216
R1767 avss.n269 avss.n268 0.00641216
R1768 avss.n281 avss.n280 0.00641216
R1769 avss.n293 avss.n292 0.00641216
R1770 avss.n304 avss.n0 0.00641216
R1771 avss.n790 avss.n354 0.004875
R1772 vin_vunder.n62 vin_vunder.t29 51.0275
R1773 vin_vunder.n7 vin_vunder.n6 48.371
R1774 vin_vunder.n20 vin_vunder.n19 48.371
R1775 vin_vunder.n14 vin_vunder.n13 48.371
R1776 vin_vunder.n10 vin_vunder.n9 48.371
R1777 vin_vunder.n74 vin_vunder.n73 48.371
R1778 vin_vunder.n70 vin_vunder.n56 48.371
R1779 vin_vunder.n67 vin_vunder.n54 48.371
R1780 vin_vunder.n77 vin_vunder.n1 48.371
R1781 vin_vunder.n22 vin_vunder.n21 45.4885
R1782 vin_vunder.n12 vin_vunder.n5 45.4885
R1783 vin_vunder.n8 vin_vunder.n4 45.4885
R1784 vin_vunder.n3 vin_vunder.n2 45.4885
R1785 vin_vunder.n55 vin_vunder.n53 45.4885
R1786 vin_vunder.n69 vin_vunder.n68 45.4885
R1787 vin_vunder.n76 vin_vunder.n75 45.4885
R1788 vin_vunder.n39 vin_vunder.n38 45.3881
R1789 vin_vunder.n63 vin_vunder.t44 20.2802
R1790 vin_vunder.n43 vin_vunder.n42 17.7666
R1791 vin_vunder.n46 vin_vunder.n45 17.7666
R1792 vin_vunder.n49 vin_vunder.n48 17.7666
R1793 vin_vunder.n59 vin_vunder.n58 17.7666
R1794 vin_vunder.n66 vin_vunder.n61 17.7666
R1795 vin_vunder.n64 vin_vunder.n63 17.7666
R1796 vin_vunder.n52 vin_vunder.n51 17.7666
R1797 vin_vunder.n39 vin_vunder.n23 17.6963
R1798 vin_vunder.n41 vin_vunder.n40 16.9742
R1799 vin_vunder.n44 vin_vunder.n43 16.9742
R1800 vin_vunder.n47 vin_vunder.n46 16.9742
R1801 vin_vunder.n50 vin_vunder.n49 16.9742
R1802 vin_vunder.n60 vin_vunder.n59 16.9742
R1803 vin_vunder.n66 vin_vunder.n65 16.9742
R1804 vin_vunder.n57 vin_vunder.n52 16.9742
R1805 vin_vunder.n31 vin_vunder.t50 9.72783
R1806 vin_vunder.n24 vin_vunder.t56 9.65028
R1807 vin_vunder.n38 vin_vunder.n30 8.96563
R1808 vin_vunder.n37 vin_vunder.t63 8.73727
R1809 vin_vunder.n36 vin_vunder.t48 8.73727
R1810 vin_vunder.n35 vin_vunder.t52 8.73727
R1811 vin_vunder.n34 vin_vunder.t60 8.73727
R1812 vin_vunder.n33 vin_vunder.t51 8.73727
R1813 vin_vunder.n32 vin_vunder.t57 8.73727
R1814 vin_vunder.n31 vin_vunder.t62 8.73727
R1815 vin_vunder.n30 vin_vunder.t54 8.65985
R1816 vin_vunder.n29 vin_vunder.t55 8.65985
R1817 vin_vunder.n28 vin_vunder.t59 8.65985
R1818 vin_vunder.n27 vin_vunder.t49 8.65985
R1819 vin_vunder.n26 vin_vunder.t58 8.65985
R1820 vin_vunder.n25 vin_vunder.t61 8.65985
R1821 vin_vunder.n24 vin_vunder.t53 8.65985
R1822 vin_vunder.n38 vin_vunder.n37 5.98511
R1823 vin_vunder.n21 vin_vunder.t43 5.5395
R1824 vin_vunder.n21 vin_vunder.t26 5.5395
R1825 vin_vunder.n6 vin_vunder.t25 5.5395
R1826 vin_vunder.n6 vin_vunder.t42 5.5395
R1827 vin_vunder.t30 vin_vunder.n12 5.5395
R1828 vin_vunder.n12 vin_vunder.t15 5.5395
R1829 vin_vunder.n20 vin_vunder.t14 5.5395
R1830 vin_vunder.t43 vin_vunder.n20 5.5395
R1831 vin_vunder.t41 vin_vunder.n8 5.5395
R1832 vin_vunder.n8 vin_vunder.t12 5.5395
R1833 vin_vunder.n13 vin_vunder.t13 5.5395
R1834 vin_vunder.n13 vin_vunder.t30 5.5395
R1835 vin_vunder.n2 vin_vunder.t27 5.5395
R1836 vin_vunder.n2 vin_vunder.t33 5.5395
R1837 vin_vunder.n9 vin_vunder.t34 5.5395
R1838 vin_vunder.n9 vin_vunder.t41 5.5395
R1839 vin_vunder.t24 vin_vunder.n55 5.5395
R1840 vin_vunder.n55 vin_vunder.t21 5.5395
R1841 vin_vunder.n74 vin_vunder.t20 5.5395
R1842 vin_vunder.t39 vin_vunder.n74 5.5395
R1843 vin_vunder.n68 vin_vunder.t40 5.5395
R1844 vin_vunder.n68 vin_vunder.t17 5.5395
R1845 vin_vunder.n56 vin_vunder.t16 5.5395
R1846 vin_vunder.n56 vin_vunder.t24 5.5395
R1847 vin_vunder.n67 vin_vunder.t28 5.5395
R1848 vin_vunder.t40 vin_vunder.n67 5.5395
R1849 vin_vunder.n75 vin_vunder.t39 5.5395
R1850 vin_vunder.n75 vin_vunder.t32 5.5395
R1851 vin_vunder.n1 vin_vunder.t31 5.5395
R1852 vin_vunder.t27 vin_vunder.n1 5.5395
R1853 vin_vunder.n71 vin_vunder.n54 3.79433
R1854 vin_vunder.n17 vin_vunder.n7 3.42225
R1855 vin_vunder.n71 vin_vunder.n70 3.4105
R1856 vin_vunder.n73 vin_vunder.n72 3.4105
R1857 vin_vunder.n78 vin_vunder.n77 3.4105
R1858 vin_vunder.n11 vin_vunder.n10 3.4105
R1859 vin_vunder.n15 vin_vunder.n14 3.4105
R1860 vin_vunder.n19 vin_vunder.n18 3.4105
R1861 vin_vunder.t1 vin_vunder.n41 3.3065
R1862 vin_vunder.n41 vin_vunder.t37 3.3065
R1863 vin_vunder.n23 vin_vunder.t38 3.3065
R1864 vin_vunder.n23 vin_vunder.t7 3.3065
R1865 vin_vunder.t3 vin_vunder.n44 3.3065
R1866 vin_vunder.n44 vin_vunder.t46 3.3065
R1867 vin_vunder.n42 vin_vunder.t47 3.3065
R1868 vin_vunder.n42 vin_vunder.t1 3.3065
R1869 vin_vunder.t5 vin_vunder.n47 3.3065
R1870 vin_vunder.n47 vin_vunder.t18 3.3065
R1871 vin_vunder.n45 vin_vunder.t19 3.3065
R1872 vin_vunder.n45 vin_vunder.t3 3.3065
R1873 vin_vunder.t2 vin_vunder.n50 3.3065
R1874 vin_vunder.n50 vin_vunder.t11 3.3065
R1875 vin_vunder.n48 vin_vunder.t10 3.3065
R1876 vin_vunder.n48 vin_vunder.t5 3.3065
R1877 vin_vunder.t4 vin_vunder.n60 3.3065
R1878 vin_vunder.n60 vin_vunder.t9 3.3065
R1879 vin_vunder.n58 vin_vunder.t8 3.3065
R1880 vin_vunder.n58 vin_vunder.t6 3.3065
R1881 vin_vunder.n65 vin_vunder.t0 3.3065
R1882 vin_vunder.n65 vin_vunder.t36 3.3065
R1883 vin_vunder.n61 vin_vunder.t35 3.3065
R1884 vin_vunder.n61 vin_vunder.t4 3.3065
R1885 vin_vunder.n64 vin_vunder.t45 3.3065
R1886 vin_vunder.t0 vin_vunder.n64 3.3065
R1887 vin_vunder.t6 vin_vunder.n57 3.3065
R1888 vin_vunder.n57 vin_vunder.t22 3.3065
R1889 vin_vunder.n51 vin_vunder.t23 3.3065
R1890 vin_vunder.n51 vin_vunder.t2 3.3065
R1891 vin_vunder.n40 vin_vunder.n22 1.98319
R1892 vin_vunder.n43 vin_vunder.n5 1.98319
R1893 vin_vunder.n46 vin_vunder.n4 1.98319
R1894 vin_vunder.n49 vin_vunder.n3 1.98319
R1895 vin_vunder.n59 vin_vunder.n53 1.98319
R1896 vin_vunder.n69 vin_vunder.n66 1.98319
R1897 vin_vunder.n63 vin_vunder.n62 1.98319
R1898 vin_vunder.n76 vin_vunder.n52 1.98319
R1899 vin_vunder.n37 vin_vunder.n36 0.99106
R1900 vin_vunder.n36 vin_vunder.n35 0.99106
R1901 vin_vunder.n35 vin_vunder.n34 0.99106
R1902 vin_vunder.n34 vin_vunder.n33 0.99106
R1903 vin_vunder.n33 vin_vunder.n32 0.99106
R1904 vin_vunder.n32 vin_vunder.n31 0.99106
R1905 vin_vunder.n30 vin_vunder.n29 0.99093
R1906 vin_vunder.n29 vin_vunder.n28 0.99093
R1907 vin_vunder.n28 vin_vunder.n27 0.99093
R1908 vin_vunder.n27 vin_vunder.n26 0.99093
R1909 vin_vunder.n26 vin_vunder.n25 0.99093
R1910 vin_vunder.n25 vin_vunder.n24 0.99093
R1911 vin_vunder.n17 vin_vunder.n16 0.678824
R1912 vin_vunder.n72 vin_vunder.n71 0.384333
R1913 vin_vunder.n15 vin_vunder.n11 0.384333
R1914 vin_vunder.n18 vin_vunder.n15 0.384333
R1915 vin_vunder.n72 vin_vunder.n0 0.372583
R1916 vin_vunder.n11 vin_vunder.n0 0.372583
R1917 vin_vunder.n18 vin_vunder.n17 0.372583
R1918 vin_vunder.n40 vin_vunder.n39 0.0708125
R1919 vin_vunder vin_vunder.n78 0.0475
R1920 vin_vunder.n78 vin_vunder.n0 0.00240541
R1921 vin_vunder.n22 vin_vunder.n7 0.00218919
R1922 vin_vunder.n19 vin_vunder.n5 0.00218919
R1923 vin_vunder.n14 vin_vunder.n4 0.00218919
R1924 vin_vunder.n10 vin_vunder.n3 0.00218919
R1925 vin_vunder.n73 vin_vunder.n53 0.00218919
R1926 vin_vunder.n70 vin_vunder.n69 0.00218919
R1927 vin_vunder.n62 vin_vunder.n54 0.00218919
R1928 vin_vunder.n77 vin_vunder.n76 0.00218919
R1929 rstring_mux_0.vtrip4.n5 rstring_mux_0.vtrip4.n3 50.7022
R1930 rstring_mux_0.vtrip4.n2 rstring_mux_0.vtrip4.n0 50.7022
R1931 rstring_mux_0.vtrip4.n7 rstring_mux_0.vtrip4.n6 24.0569
R1932 rstring_mux_0.vtrip4.n6 rstring_mux_0.vtrip4.n2 14.0584
R1933 rstring_mux_0.vtrip4.n5 rstring_mux_0.vtrip4.n4 13.8791
R1934 rstring_mux_0.vtrip4.n2 rstring_mux_0.vtrip4.n1 13.8791
R1935 rstring_mux_0.vtrip4.n7 rstring_mux_0.vtrip4.t9 10.6303
R1936 rstring_mux_0.vtrip4.n3 rstring_mux_0.vtrip4.t1 5.5395
R1937 rstring_mux_0.vtrip4.n3 rstring_mux_0.vtrip4.t2 5.5395
R1938 rstring_mux_0.vtrip4.n0 rstring_mux_0.vtrip4.t6 5.5395
R1939 rstring_mux_0.vtrip4.n0 rstring_mux_0.vtrip4.t5 5.5395
R1940 rstring_mux_0.vtrip4.n6 rstring_mux_0.vtrip4.n5 3.33746
R1941 rstring_mux_0.vtrip4.n4 rstring_mux_0.vtrip4.t8 3.3065
R1942 rstring_mux_0.vtrip4.n4 rstring_mux_0.vtrip4.t7 3.3065
R1943 rstring_mux_0.vtrip4.n1 rstring_mux_0.vtrip4.t3 3.3065
R1944 rstring_mux_0.vtrip4.n1 rstring_mux_0.vtrip4.t4 3.3065
R1945 rstring_mux_0.vtrip4 rstring_mux_0.vtrip4.t0 0.769662
R1946 rstring_mux_0.vtrip4 rstring_mux_0.vtrip4.n7 0.0563195
R1947 avdd.n1494 avdd.n1450 99969.2
R1948 avdd.n1494 avdd.n1493 83663.1
R1949 avdd.n1478 avdd.n1451 66867
R1950 avdd.n1479 avdd.n1452 60783.5
R1951 avdd.n1478 avdd.n1477 60384.8
R1952 avdd.n1467 avdd.n1450 58787
R1953 avdd.n1491 avdd.n1452 52810.3
R1954 avdd.n1492 avdd.n1451 50831
R1955 avdd.n1495 avdd.n1448 49200
R1956 avdd.n1477 avdd.n1476 47131.3
R1957 avdd.n1495 avdd.n1449 41239.5
R1958 avdd.n1479 avdd.n1457 29875.1
R1959 avdd.n1468 avdd.n1448 29132.4
R1960 avdd.n1493 avdd.n1492 27601.7
R1961 avdd.n1467 avdd.n1458 27058.6
R1962 avdd.n1144 avdd.n1017 25108.6
R1963 avdd.n1142 avdd.n1017 25108.6
R1964 avdd.n1390 avdd.n1263 25108.6
R1965 avdd.n1388 avdd.n1263 25108.6
R1966 avdd.n1144 avdd.n1143 25105.2
R1967 avdd.n1143 avdd.n1142 25105.2
R1968 avdd.n1390 avdd.n1389 25105.2
R1969 avdd.n1389 avdd.n1388 25105.2
R1970 avdd.n1475 avdd.n1457 22957.3
R1971 avdd.n1476 avdd.n1458 17438.8
R1972 avdd.n1546 avdd.n1539 15077.5
R1973 avdd.n1546 avdd.n1540 15077.5
R1974 avdd.n1583 avdd.n1540 15077.5
R1975 avdd.n1583 avdd.n1539 15077.5
R1976 avdd.n1491 avdd.n1449 13877.8
R1977 avdd.n1468 avdd.n1459 13642.7
R1978 avdd.n1145 avdd.n1015 12653.5
R1979 avdd.n1141 avdd.n1015 12653.5
R1980 avdd.n1391 avdd.n1261 12653.5
R1981 avdd.n1387 avdd.n1261 12653.5
R1982 avdd.n1145 avdd.n1016 12651.9
R1983 avdd.n1141 avdd.n1016 12651.9
R1984 avdd.n1391 avdd.n1262 12651.9
R1985 avdd.n1387 avdd.n1262 12651.9
R1986 avdd.n1165 avdd.n962 11582.8
R1987 avdd.n1125 avdd.n962 11582.8
R1988 avdd.n1411 avdd.n1208 11582.8
R1989 avdd.n1371 avdd.n1208 11582.8
R1990 avdd.n1167 avdd.n959 10507.7
R1991 avdd.n1127 avdd.n959 10507.7
R1992 avdd.n1413 avdd.n1205 10507.7
R1993 avdd.n1373 avdd.n1205 10507.7
R1994 avdd.n1159 avdd.n979 10039.9
R1995 avdd.n1159 avdd.n958 10039.9
R1996 avdd.n1161 avdd.n978 10039.9
R1997 avdd.n1161 avdd.n963 10039.9
R1998 avdd.n1405 avdd.n1225 10039.9
R1999 avdd.n1405 avdd.n1204 10039.9
R2000 avdd.n1407 avdd.n1224 10039.9
R2001 avdd.n1407 avdd.n1209 10039.9
R2002 avdd.n1647 avdd.n692 9739.14
R2003 avdd.n1647 avdd.n693 9739.14
R2004 avdd.n1646 avdd.n693 9739.14
R2005 avdd.n1646 avdd.n692 9739.14
R2006 avdd.n1475 avdd.n1459 8461.62
R2007 avdd.n1481 avdd.n1453 8070.02
R2008 avdd.n1480 avdd.n1456 6943.25
R2009 avdd.n1466 avdd.n1465 6761.04
R2010 avdd.n1490 avdd.n1453 6168.09
R2011 avdd.n1473 avdd.n1461 5303.72
R2012 avdd.n1486 avdd.n1485 4892.23
R2013 avdd.n1497 avdd.n1446 4681.79
R2014 avdd.n1463 avdd.n1446 4335.44
R2015 avdd.n1631 avdd.n1630 4316.28
R2016 avdd.n1633 avdd.n1630 4316.28
R2017 avdd.n1631 avdd.n1627 4316.28
R2018 avdd.n1633 avdd.n1627 4316.28
R2019 avdd.n1489 avdd.n1454 3225.22
R2020 avdd.n1470 avdd.n1469 3163.48
R2021 avdd.n1598 avdd.n1511 3160.55
R2022 avdd.n1599 avdd.n1511 3160.55
R2023 avdd.n1146 avdd.n1014 2933.46
R2024 avdd.n1392 avdd.n1260 2933.46
R2025 avdd.n1140 avdd.n1018 2922.54
R2026 avdd.n1386 avdd.n1264 2922.54
R2027 avdd.n1582 avdd.n1541 2890.84
R2028 avdd.n1547 avdd.n1541 2890.84
R2029 avdd.n1139 avdd.n1019 2865.69
R2030 avdd.n1385 avdd.n1265 2865.69
R2031 avdd.n1548 avdd.n1542 2860.42
R2032 avdd.n1581 avdd.n1542 2860.42
R2033 avdd.n1147 avdd.n1013 2841.22
R2034 avdd.n1393 avdd.n1259 2841.22
R2035 avdd.n1123 avdd.n978 2620.03
R2036 avdd.n1123 avdd.n979 2620.03
R2037 avdd.n963 avdd.n960 2620.03
R2038 avdd.n960 avdd.n958 2620.03
R2039 avdd.n1369 avdd.n1224 2620.03
R2040 avdd.n1369 avdd.n1225 2620.03
R2041 avdd.n1209 avdd.n1206 2620.03
R2042 avdd.n1206 avdd.n1204 2620.03
R2043 avdd.n1592 avdd.n1518 2513.9
R2044 avdd.n1592 avdd.n1510 2513.9
R2045 avdd.n1593 avdd.n1515 2513.9
R2046 avdd.n1593 avdd.n1512 2513.9
R2047 avdd.n1485 avdd.n1447 2495.62
R2048 avdd.n1121 avdd.n1036 2480.48
R2049 avdd.n1121 avdd.n1037 2480.48
R2050 avdd.n1036 avdd.n1035 2480.48
R2051 avdd.n1037 avdd.n1035 2480.48
R2052 avdd.n1367 avdd.n1282 2480.48
R2053 avdd.n1367 avdd.n1283 2480.48
R2054 avdd.n1282 avdd.n1281 2480.48
R2055 avdd.n1283 avdd.n1281 2480.48
R2056 avdd.n1497 avdd.n1496 2412.42
R2057 avdd.n1587 avdd.n1535 2346.83
R2058 avdd.n1586 avdd.n1535 2346.83
R2059 avdd.n1124 avdd.n964 2223.06
R2060 avdd.n1164 avdd.n964 2223.06
R2061 avdd.n1370 avdd.n1210 2223.06
R2062 avdd.n1410 avdd.n1210 2223.06
R2063 avdd.n1496 avdd.n1447 2115.76
R2064 avdd.n972 avdd.n971 2059.86
R2065 avdd.n971 avdd.n970 2059.86
R2066 avdd.n970 avdd.n967 2059.86
R2067 avdd.n972 avdd.n967 2059.86
R2068 avdd.n1218 avdd.n1217 2059.86
R2069 avdd.n1217 avdd.n1216 2059.86
R2070 avdd.n1216 avdd.n1213 2059.86
R2071 avdd.n1218 avdd.n1213 2059.86
R2072 avdd.n1168 avdd.n957 2000.19
R2073 avdd.n1128 avdd.n957 2000.19
R2074 avdd.n1414 avdd.n1203 2000.19
R2075 avdd.n1374 avdd.n1203 2000.19
R2076 avdd.n1474 avdd.n1460 1971.95
R2077 avdd.n1162 avdd.n976 1923.01
R2078 avdd.n1163 avdd.n1162 1923.01
R2079 avdd.n1408 avdd.n1222 1923.01
R2080 avdd.n1409 avdd.n1408 1923.01
R2081 avdd.n1599 avdd.n1510 1837.76
R2082 avdd.n1598 avdd.n1512 1837.76
R2083 avdd.n694 avdd.n690 1616.56
R2084 avdd.n1644 avdd.n695 1616.56
R2085 avdd.n695 avdd.n691 1616.56
R2086 avdd.n1649 avdd.n690 1615.06
R2087 avdd.n1165 avdd.n963 1542.93
R2088 avdd.n1125 avdd.n978 1542.93
R2089 avdd.n1411 avdd.n1209 1542.93
R2090 avdd.n1371 avdd.n1224 1542.93
R2091 avdd.n1537 avdd.n1515 1322.79
R2092 avdd.n1537 avdd.n1518 1322.79
R2093 avdd.n1516 avdd.n1512 1322.79
R2094 avdd.n1516 avdd.n1510 1322.79
R2095 avdd.n1158 avdd.n980 1237.08
R2096 avdd.n1158 avdd.n955 1237.08
R2097 avdd.n1404 avdd.n1226 1237.08
R2098 avdd.n1404 avdd.n1201 1237.08
R2099 avdd.n1587 avdd.n1518 1024.03
R2100 avdd.n1586 avdd.n1515 1024.03
R2101 avdd.n1635 avdd.n1634 831.247
R2102 avdd.n1635 avdd.n1626 831.247
R2103 avdd.n73 avdd.t166 692.692
R2104 avdd.n409 avdd.t162 692.692
R2105 avdd avdd.t169 688.231
R2106 avdd avdd.t49 688.231
R2107 avdd.n1629 avdd.n1628 682.918
R2108 avdd.n1629 avdd.n1609 682.918
R2109 avdd.n334 avdd.t160 648.668
R2110 avdd.n306 avdd.t520 648.668
R2111 avdd.n278 avdd.t453 648.668
R2112 avdd.n250 avdd.t585 648.668
R2113 avdd.n222 avdd.t405 648.668
R2114 avdd.n194 avdd.t121 648.668
R2115 avdd.n166 avdd.t514 648.668
R2116 avdd.n138 avdd.t487 648.668
R2117 avdd.n110 avdd.t51 648.668
R2118 avdd.n670 avdd.t417 648.668
R2119 avdd.n642 avdd.t497 648.668
R2120 avdd.n614 avdd.t441 648.668
R2121 avdd.n586 avdd.t536 648.668
R2122 avdd.n558 avdd.t115 648.668
R2123 avdd.n530 avdd.t57 648.668
R2124 avdd.n502 avdd.t608 648.668
R2125 avdd.n474 avdd.t13 648.668
R2126 avdd.n446 avdd.t7 648.668
R2127 avdd.n922 avdd.n705 624.808
R2128 avdd.n920 avdd.n706 624.808
R2129 avdd.n909 avdd.n908 624.808
R2130 avdd.n897 avdd.n725 624.808
R2131 avdd.n895 avdd.n726 624.808
R2132 avdd.n884 avdd.n883 624.808
R2133 avdd.n872 avdd.n745 624.808
R2134 avdd.n870 avdd.n746 624.808
R2135 avdd.n859 avdd.n858 624.808
R2136 avdd.n847 avdd.n765 624.808
R2137 avdd.n845 avdd.n766 624.808
R2138 avdd.n834 avdd.n833 624.808
R2139 avdd.n822 avdd.n785 624.808
R2140 avdd.n820 avdd.n786 624.808
R2141 avdd.n809 avdd.n808 624.808
R2142 avdd.n1130 avdd.n980 612.894
R2143 avdd.n1170 avdd.n955 612.894
R2144 avdd.n1376 avdd.n1226 612.894
R2145 avdd.n1416 avdd.n1201 612.894
R2146 avdd.n1597 avdd.n1508 609.883
R2147 avdd.n1601 avdd.n1600 555.672
R2148 avdd.t92 avdd.t90 511.356
R2149 avdd.t336 avdd.t98 511.356
R2150 avdd.t505 avdd.t336 511.356
R2151 avdd.t507 avdd.t505 511.356
R2152 avdd.t371 avdd.t507 511.356
R2153 avdd.t509 avdd.t371 511.356
R2154 avdd.t511 avdd.t509 511.356
R2155 avdd.t264 avdd.t511 511.356
R2156 avdd.n1129 avdd.n1034 506.353
R2157 avdd.n1375 avdd.n1280 506.353
R2158 avdd.n680 avdd.t541 499.882
R2159 avdd.t543 avdd.t551 484.288
R2160 avdd.t174 avdd.t549 484.288
R2161 avdd.t561 avdd.t553 484.288
R2162 avdd.t524 avdd.t559 484.288
R2163 avdd.n1591 avdd.n1589 481.507
R2164 avdd.n1594 avdd.n1514 481.507
R2165 avdd.n1041 avdd.n1040 479.625
R2166 avdd.n1040 avdd.n1039 479.625
R2167 avdd.n1287 avdd.n1286 479.625
R2168 avdd.n1286 avdd.n1285 479.625
R2169 avdd.t90 avdd.t94 475.098
R2170 avdd.n1167 avdd.n958 467.793
R2171 avdd.n1127 avdd.n979 467.793
R2172 avdd.n1413 avdd.n1204 467.793
R2173 avdd.n1373 avdd.n1225 467.793
R2174 avdd.n1585 avdd.n1534 454.024
R2175 avdd.n970 avdd.t174 437.699
R2176 avdd.n1216 avdd.t524 437.699
R2177 avdd.n1120 avdd.n1038 437.082
R2178 avdd.n1120 avdd.n1119 437.082
R2179 avdd.n1366 avdd.n1284 437.082
R2180 avdd.n1366 avdd.n1365 437.082
R2181 avdd.n1588 avdd.n1534 423.818
R2182 avdd.n973 avdd.n966 399.06
R2183 avdd.n969 avdd.n966 399.06
R2184 avdd.n1219 avdd.n1212 399.06
R2185 avdd.n1215 avdd.n1212 399.06
R2186 avdd.n1522 avdd.t343 397.264
R2187 avdd.n1523 avdd.t350 397.135
R2188 avdd.n1524 avdd.t233 397.135
R2189 avdd.n689 avdd.t253 388.149
R2190 avdd.n933 avdd.t362 388.149
R2191 avdd.n934 avdd.t400 388.149
R2192 avdd.n935 avdd.t396 388.149
R2193 avdd.n936 avdd.t302 388.149
R2194 avdd.n937 avdd.t384 388.149
R2195 avdd.n938 avdd.t373 388.149
R2196 avdd.n939 avdd.t386 388.149
R2197 avdd.n941 avdd.t398 388.149
R2198 avdd.n942 avdd.t267 388.149
R2199 avdd.n943 avdd.t380 388.149
R2200 avdd.n944 avdd.t280 388.149
R2201 avdd.n945 avdd.t338 388.149
R2202 avdd.n946 avdd.t248 388.149
R2203 avdd.n947 avdd.t309 388.149
R2204 avdd.n330 avdd.t15 372.885
R2205 avdd.n302 avdd.t457 372.885
R2206 avdd.n274 avdd.t210 372.885
R2207 avdd.n246 avdd.t445 372.885
R2208 avdd.n218 avdd.t485 372.885
R2209 avdd.n190 avdd.t206 372.885
R2210 avdd.n162 avdd.t415 372.885
R2211 avdd.n134 avdd.t502 372.885
R2212 avdd.n106 avdd.t422 372.885
R2213 avdd.n666 avdd.t17 372.885
R2214 avdd.n638 avdd.t483 372.885
R2215 avdd.n610 avdd.t411 372.885
R2216 avdd.n582 avdd.t494 372.885
R2217 avdd.n554 avdd.t5 372.885
R2218 avdd.n526 avdd.t568 372.885
R2219 avdd.n498 avdd.t225 372.885
R2220 avdd.n470 avdd.t527 372.885
R2221 avdd.n442 avdd.t103 372.885
R2222 avdd.t563 avdd.n697 354.904
R2223 avdd.n1600 avdd.n1509 352
R2224 avdd.n1597 avdd.n1596 352
R2225 avdd.n1546 avdd.t264 345.817
R2226 avdd.n972 avdd.t543 343.495
R2227 avdd.n1218 avdd.t561 343.495
R2228 avdd.n1590 avdd.n1509 325.647
R2229 avdd.n1596 avdd.n1595 325.647
R2230 avdd.n1036 avdd.t430 323.445
R2231 avdd.n1037 avdd.t175 323.445
R2232 avdd.n1282 avdd.t592 323.445
R2233 avdd.n1283 avdd.t602 323.445
R2234 avdd.n323 avdd.n6 321.882
R2235 avdd.n309 avdd.n308 321.882
R2236 avdd.n4 avdd.n2 321.882
R2237 avdd.n295 avdd.n14 321.882
R2238 avdd.n281 avdd.n280 321.882
R2239 avdd.n12 avdd.n10 321.882
R2240 avdd.n267 avdd.n22 321.882
R2241 avdd.n253 avdd.n252 321.882
R2242 avdd.n20 avdd.n18 321.882
R2243 avdd.n239 avdd.n30 321.882
R2244 avdd.n225 avdd.n224 321.882
R2245 avdd.n28 avdd.n26 321.882
R2246 avdd.n211 avdd.n38 321.882
R2247 avdd.n197 avdd.n196 321.882
R2248 avdd.n36 avdd.n34 321.882
R2249 avdd.n183 avdd.n46 321.882
R2250 avdd.n169 avdd.n168 321.882
R2251 avdd.n44 avdd.n42 321.882
R2252 avdd.n155 avdd.n54 321.882
R2253 avdd.n141 avdd.n140 321.882
R2254 avdd.n52 avdd.n50 321.882
R2255 avdd.n127 avdd.n62 321.882
R2256 avdd.n113 avdd.n112 321.882
R2257 avdd.n60 avdd.n58 321.882
R2258 avdd.n75 avdd.n70 321.882
R2259 avdd.n92 avdd.n70 321.882
R2260 avdd.n92 avdd.n67 321.882
R2261 avdd.n96 avdd.n67 321.882
R2262 avdd.n97 avdd.n96 321.882
R2263 avdd.n97 avdd.n66 321.882
R2264 avdd.n101 avdd.n66 321.882
R2265 avdd.n659 avdd.n342 321.882
R2266 avdd.n645 avdd.n644 321.882
R2267 avdd.n340 avdd.n338 321.882
R2268 avdd.n631 avdd.n350 321.882
R2269 avdd.n617 avdd.n616 321.882
R2270 avdd.n348 avdd.n346 321.882
R2271 avdd.n603 avdd.n358 321.882
R2272 avdd.n589 avdd.n588 321.882
R2273 avdd.n356 avdd.n354 321.882
R2274 avdd.n575 avdd.n366 321.882
R2275 avdd.n561 avdd.n560 321.882
R2276 avdd.n364 avdd.n362 321.882
R2277 avdd.n547 avdd.n374 321.882
R2278 avdd.n533 avdd.n532 321.882
R2279 avdd.n372 avdd.n370 321.882
R2280 avdd.n519 avdd.n382 321.882
R2281 avdd.n505 avdd.n504 321.882
R2282 avdd.n380 avdd.n378 321.882
R2283 avdd.n491 avdd.n390 321.882
R2284 avdd.n477 avdd.n476 321.882
R2285 avdd.n388 avdd.n386 321.882
R2286 avdd.n463 avdd.n398 321.882
R2287 avdd.n449 avdd.n448 321.882
R2288 avdd.n396 avdd.n394 321.882
R2289 avdd.n411 avdd.n406 321.882
R2290 avdd.n428 avdd.n403 321.882
R2291 avdd.n432 avdd.n403 321.882
R2292 avdd.n433 avdd.n432 321.882
R2293 avdd.n433 avdd.n402 321.882
R2294 avdd.n437 avdd.n402 321.882
R2295 avdd.n679 avdd.n678 321.882
R2296 avdd.n807 avdd.n791 321.882
R2297 avdd.n812 avdd.n811 321.882
R2298 avdd.n811 avdd.n790 321.882
R2299 avdd.n823 avdd.n782 321.882
R2300 avdd.n819 avdd.n782 321.882
R2301 avdd.n832 avdd.n771 321.882
R2302 avdd.n784 avdd.n771 321.882
R2303 avdd.n837 avdd.n836 321.882
R2304 avdd.n836 avdd.n770 321.882
R2305 avdd.n848 avdd.n762 321.882
R2306 avdd.n844 avdd.n762 321.882
R2307 avdd.n857 avdd.n751 321.882
R2308 avdd.n764 avdd.n751 321.882
R2309 avdd.n862 avdd.n861 321.882
R2310 avdd.n861 avdd.n750 321.882
R2311 avdd.n873 avdd.n742 321.882
R2312 avdd.n869 avdd.n742 321.882
R2313 avdd.n882 avdd.n731 321.882
R2314 avdd.n744 avdd.n731 321.882
R2315 avdd.n887 avdd.n886 321.882
R2316 avdd.n886 avdd.n730 321.882
R2317 avdd.n898 avdd.n722 321.882
R2318 avdd.n894 avdd.n722 321.882
R2319 avdd.n907 avdd.n711 321.882
R2320 avdd.n724 avdd.n711 321.882
R2321 avdd.n912 avdd.n911 321.882
R2322 avdd.n911 avdd.n710 321.882
R2323 avdd.n923 avdd.n703 321.882
R2324 avdd.n919 avdd.n703 321.882
R2325 avdd.n698 avdd.n697 321.882
R2326 avdd.n699 avdd.n698 321.882
R2327 avdd.n799 avdd.n798 318.757
R2328 avdd.n428 avdd.n406 318.529
R2329 avdd.t246 avdd.t25 310.303
R2330 avdd.t25 avdd.t22 310.303
R2331 avdd.t18 avdd.t33 310.303
R2332 avdd.t33 avdd.t227 310.303
R2333 avdd.t240 avdd.t140 310.303
R2334 avdd.t140 avdd.t133 310.303
R2335 avdd.t125 avdd.t123 310.303
R2336 avdd.t123 avdd.t236 310.303
R2337 avdd.n1124 avdd.n976 300.048
R2338 avdd.n1164 avdd.n1163 300.048
R2339 avdd.n974 avdd.n965 300.048
R2340 avdd.n968 avdd.n965 300.048
R2341 avdd.n1370 avdd.n1222 300.048
R2342 avdd.n1410 avdd.n1409 300.048
R2343 avdd.n1220 avdd.n1211 300.048
R2344 avdd.n1214 avdd.n1211 300.048
R2345 avdd.n1033 avdd.n976 295.529
R2346 avdd.n1279 avdd.n1222 295.529
R2347 avdd.t551 avdd.n961 289.247
R2348 avdd.t553 avdd.n1207 289.247
R2349 avdd.n1169 avdd.n956 281.601
R2350 avdd.n1415 avdd.n1202 281.601
R2351 avdd.n326 avdd.n325 271.068
R2352 avdd.n298 avdd.n297 271.068
R2353 avdd.n270 avdd.n269 271.068
R2354 avdd.n242 avdd.n241 271.068
R2355 avdd.n214 avdd.n213 271.068
R2356 avdd.n186 avdd.n185 271.068
R2357 avdd.n158 avdd.n157 271.068
R2358 avdd.n130 avdd.n129 271.068
R2359 avdd.n662 avdd.n661 271.068
R2360 avdd.n634 avdd.n633 271.068
R2361 avdd.n606 avdd.n605 271.068
R2362 avdd.n578 avdd.n577 271.068
R2363 avdd.n550 avdd.n549 271.068
R2364 avdd.n522 avdd.n521 271.068
R2365 avdd.n494 avdd.n493 271.068
R2366 avdd.n466 avdd.n465 271.068
R2367 avdd.n682 avdd.n681 271.068
R2368 avdd.n1596 avdd.n1513 257.882
R2369 avdd.n1536 avdd.n1514 257.882
R2370 avdd.n1545 avdd.t92 255.679
R2371 avdd.t98 avdd.n1545 255.679
R2372 avdd.n686 avdd.t542 252.983
R2373 avdd.n802 avdd.t533 252.983
R2374 avdd.n795 avdd.t212 252.983
R2375 avdd.n815 avdd.t107 252.983
R2376 avdd.n827 avdd.t582 252.983
R2377 avdd.n775 avdd.t580 252.983
R2378 avdd.n840 avdd.t119 252.983
R2379 avdd.n852 avdd.t208 252.983
R2380 avdd.n755 avdd.t610 252.983
R2381 avdd.n865 avdd.t540 252.983
R2382 avdd.n877 avdd.t578 252.983
R2383 avdd.n735 avdd.t158 252.983
R2384 avdd.n890 avdd.t105 252.983
R2385 avdd.n902 avdd.t409 252.983
R2386 avdd.n715 avdd.t47 252.983
R2387 avdd.n915 avdd.t531 252.983
R2388 avdd.n926 avdd.t564 252.983
R2389 avdd.n1649 avdd.n1648 241.459
R2390 avdd.n1645 avdd.n694 240.66
R2391 avdd.n1645 avdd.n1644 240.66
R2392 avdd.n1648 avdd.n691 240.66
R2393 avdd.t430 avdd.t424 233.565
R2394 avdd.t424 avdd.t434 233.565
R2395 avdd.t434 avdd.t432 233.565
R2396 avdd.t432 avdd.t426 233.565
R2397 avdd.t428 avdd.t436 233.565
R2398 avdd.t438 avdd.t428 233.565
R2399 avdd.t177 avdd.t438 233.565
R2400 avdd.t175 avdd.t177 233.565
R2401 avdd.t592 avdd.t596 233.565
R2402 avdd.t596 avdd.t600 233.565
R2403 avdd.t600 avdd.t586 233.565
R2404 avdd.t586 avdd.t590 233.565
R2405 avdd.t588 avdd.t598 233.565
R2406 avdd.t594 avdd.t588 233.565
R2407 avdd.t604 avdd.t594 233.565
R2408 avdd.t602 avdd.t604 233.565
R2409 avdd.n1195 avdd.t550 232.686
R2410 avdd.n1441 avdd.t560 232.686
R2411 avdd.n1109 avdd.t431 231.989
R2412 avdd.n1118 avdd.t176 231.989
R2413 avdd.n1355 avdd.t593 231.989
R2414 avdd.n1364 avdd.t603 231.989
R2415 avdd.n1196 avdd.t544 231.974
R2416 avdd.n1195 avdd.t552 231.974
R2417 avdd.n1442 avdd.t562 231.974
R2418 avdd.n1441 avdd.t554 231.974
R2419 avdd.n1192 avdd.t252 227.478
R2420 avdd.n1190 avdd.t262 227.478
R2421 avdd.n1188 avdd.t259 227.478
R2422 avdd.n1186 avdd.t296 227.478
R2423 avdd.n1184 avdd.t316 227.478
R2424 avdd.n1182 avdd.t319 227.478
R2425 avdd.n1180 avdd.t334 227.478
R2426 avdd.n1178 avdd.t329 227.478
R2427 avdd.n1176 avdd.t390 227.478
R2428 avdd.n1174 avdd.t342 227.478
R2429 avdd.n1172 avdd.t395 227.478
R2430 avdd.n1105 avdd.t283 227.478
R2431 avdd.t290 avdd.n1100 227.478
R2432 avdd.t288 avdd.n1097 227.478
R2433 avdd.n1094 avdd.t353 227.478
R2434 avdd.n1091 avdd.t367 227.478
R2435 avdd.t369 avdd.n1086 227.478
R2436 avdd.t383 avdd.n1083 227.478
R2437 avdd.n1080 avdd.t376 227.478
R2438 avdd.n1077 avdd.t247 227.478
R2439 avdd.t392 avdd.n1072 227.478
R2440 avdd.t256 avdd.n1069 227.478
R2441 avdd.n1438 avdd.t322 227.478
R2442 avdd.n1436 avdd.t299 227.478
R2443 avdd.n1434 avdd.t313 227.478
R2444 avdd.n1432 avdd.t293 227.478
R2445 avdd.n1430 avdd.t244 227.478
R2446 avdd.n1428 avdd.t286 227.478
R2447 avdd.n1426 avdd.t238 227.478
R2448 avdd.n1424 avdd.t379 227.478
R2449 avdd.n1422 avdd.t361 227.478
R2450 avdd.n1420 avdd.t358 227.478
R2451 avdd.n1418 avdd.t306 227.478
R2452 avdd.n1351 avdd.t365 227.478
R2453 avdd.t349 avdd.n1346 227.478
R2454 avdd.t355 avdd.n1343 227.478
R2455 avdd.n1340 avdd.t347 227.478
R2456 avdd.n1337 avdd.t276 227.478
R2457 avdd.t331 avdd.n1332 227.478
R2458 avdd.t272 avdd.n1329 227.478
R2459 avdd.n1326 avdd.t326 227.478
R2460 avdd.n1323 avdd.t308 227.478
R2461 avdd.t301 avdd.n1318 227.478
R2462 avdd.t270 avdd.n1315 227.478
R2463 avdd.n953 avdd.t229 227.345
R2464 avdd.t274 avdd.n1133 227.345
R2465 avdd.n1199 avdd.t279 227.345
R2466 avdd.t241 avdd.n1379 227.345
R2467 avdd.n1026 avdd.n956 211.953
R2468 avdd.n1272 avdd.n1202 211.953
R2469 avdd.n1588 avdd.t323 211.924
R2470 avdd.n1034 avdd.n1033 210.825
R2471 avdd.n1280 avdd.n1279 210.825
R2472 avdd.n1156 avdd.n1155 204.31
R2473 avdd.n1135 avdd.n1134 204.31
R2474 avdd.n1010 avdd.n1009 204.31
R2475 avdd.n1402 avdd.n1401 204.31
R2476 avdd.n1381 avdd.n1380 204.31
R2477 avdd.n1256 avdd.n1255 204.31
R2478 avdd.n1111 avdd.n1110 204.294
R2479 avdd.n1113 avdd.n1112 204.294
R2480 avdd.n1115 avdd.n1114 204.294
R2481 avdd.n1117 avdd.n1116 204.294
R2482 avdd.n1357 avdd.n1356 204.294
R2483 avdd.n1359 avdd.n1358 204.294
R2484 avdd.n1361 avdd.n1360 204.294
R2485 avdd.n1363 avdd.n1362 204.294
R2486 avdd.n1061 avdd.n1060 204.284
R2487 avdd.n1059 avdd.n1058 204.284
R2488 avdd.n1057 avdd.n1056 204.284
R2489 avdd.n1055 avdd.n1054 204.284
R2490 avdd.n1053 avdd.n1052 204.284
R2491 avdd.n1051 avdd.n1050 204.284
R2492 avdd.n1049 avdd.n1048 204.284
R2493 avdd.n1047 avdd.n1046 204.284
R2494 avdd.n1045 avdd.n1044 204.284
R2495 avdd.n1043 avdd.n1042 204.284
R2496 avdd.n982 avdd.n981 204.284
R2497 avdd.n1104 avdd.n1103 204.284
R2498 avdd.n1102 avdd.n1101 204.284
R2499 avdd.n1099 avdd.n1098 204.284
R2500 avdd.n1093 avdd.n1065 204.284
R2501 avdd.n1090 avdd.n1089 204.284
R2502 avdd.n1088 avdd.n1087 204.284
R2503 avdd.n1085 avdd.n1084 204.284
R2504 avdd.n1079 avdd.n1067 204.284
R2505 avdd.n1076 avdd.n1075 204.284
R2506 avdd.n1074 avdd.n1073 204.284
R2507 avdd.n1071 avdd.n1070 204.284
R2508 avdd.n987 avdd.n986 204.284
R2509 avdd.n989 avdd.n988 204.284
R2510 avdd.n991 avdd.n990 204.284
R2511 avdd.n993 avdd.n992 204.284
R2512 avdd.n995 avdd.n994 204.284
R2513 avdd.n997 avdd.n996 204.284
R2514 avdd.n999 avdd.n998 204.284
R2515 avdd.n1001 avdd.n1000 204.284
R2516 avdd.n1003 avdd.n1002 204.284
R2517 avdd.n1005 avdd.n1004 204.284
R2518 avdd.n1007 avdd.n1006 204.284
R2519 avdd.n1307 avdd.n1306 204.284
R2520 avdd.n1305 avdd.n1304 204.284
R2521 avdd.n1303 avdd.n1302 204.284
R2522 avdd.n1301 avdd.n1300 204.284
R2523 avdd.n1299 avdd.n1298 204.284
R2524 avdd.n1297 avdd.n1296 204.284
R2525 avdd.n1295 avdd.n1294 204.284
R2526 avdd.n1293 avdd.n1292 204.284
R2527 avdd.n1291 avdd.n1290 204.284
R2528 avdd.n1289 avdd.n1288 204.284
R2529 avdd.n1228 avdd.n1227 204.284
R2530 avdd.n1350 avdd.n1349 204.284
R2531 avdd.n1348 avdd.n1347 204.284
R2532 avdd.n1345 avdd.n1344 204.284
R2533 avdd.n1339 avdd.n1311 204.284
R2534 avdd.n1336 avdd.n1335 204.284
R2535 avdd.n1334 avdd.n1333 204.284
R2536 avdd.n1331 avdd.n1330 204.284
R2537 avdd.n1325 avdd.n1313 204.284
R2538 avdd.n1322 avdd.n1321 204.284
R2539 avdd.n1320 avdd.n1319 204.284
R2540 avdd.n1317 avdd.n1316 204.284
R2541 avdd.n1233 avdd.n1232 204.284
R2542 avdd.n1235 avdd.n1234 204.284
R2543 avdd.n1237 avdd.n1236 204.284
R2544 avdd.n1239 avdd.n1238 204.284
R2545 avdd.n1241 avdd.n1240 204.284
R2546 avdd.n1243 avdd.n1242 204.284
R2547 avdd.n1245 avdd.n1244 204.284
R2548 avdd.n1247 avdd.n1246 204.284
R2549 avdd.n1249 avdd.n1248 204.284
R2550 avdd.n1251 avdd.n1250 204.284
R2551 avdd.n1253 avdd.n1252 204.284
R2552 avdd.n1525 avdd.n1509 203.672
R2553 avdd.n1589 avdd.n1533 203.672
R2554 avdd.n1027 avdd.n1026 201.788
R2555 avdd.n1273 avdd.n1272 201.788
R2556 avdd.n324 avdd.t14 197.562
R2557 avdd.n296 avdd.t456 197.562
R2558 avdd.n268 avdd.t209 197.562
R2559 avdd.n240 avdd.t444 197.562
R2560 avdd.n212 avdd.t484 197.562
R2561 avdd.n184 avdd.t205 197.562
R2562 avdd.n156 avdd.t414 197.562
R2563 avdd.n128 avdd.t501 197.562
R2564 avdd.n660 avdd.t16 197.562
R2565 avdd.n632 avdd.t482 197.562
R2566 avdd.n604 avdd.t410 197.562
R2567 avdd.n576 avdd.t493 197.562
R2568 avdd.n548 avdd.t4 197.562
R2569 avdd.n520 avdd.t567 197.562
R2570 avdd.n492 avdd.t224 197.562
R2571 avdd.n464 avdd.t526 197.562
R2572 avdd.n1585 avdd.n1514 196.142
R2573 avdd.t549 avdd.n961 195.042
R2574 avdd.t559 avdd.n1207 195.042
R2575 avdd.n75 avdd.t165 193.774
R2576 avdd.n411 avdd.t48 193.774
R2577 avdd.n1027 avdd.n975 186.353
R2578 avdd.n1273 avdd.n1221 186.353
R2579 avdd.n323 avdd.n322 185
R2580 avdd.n324 avdd.n323 185
R2581 avdd.n7 avdd.n6 185
R2582 avdd.n318 avdd.n308 185
R2583 avdd.n317 avdd.n309 185
R2584 avdd.n4 avdd.n1 185
R2585 avdd.n327 avdd.n2 185
R2586 avdd.n295 avdd.n294 185
R2587 avdd.n296 avdd.n295 185
R2588 avdd.n15 avdd.n14 185
R2589 avdd.n290 avdd.n280 185
R2590 avdd.n289 avdd.n281 185
R2591 avdd.n12 avdd.n9 185
R2592 avdd.n299 avdd.n10 185
R2593 avdd.n267 avdd.n266 185
R2594 avdd.n268 avdd.n267 185
R2595 avdd.n23 avdd.n22 185
R2596 avdd.n262 avdd.n252 185
R2597 avdd.n261 avdd.n253 185
R2598 avdd.n20 avdd.n17 185
R2599 avdd.n271 avdd.n18 185
R2600 avdd.n239 avdd.n238 185
R2601 avdd.n240 avdd.n239 185
R2602 avdd.n31 avdd.n30 185
R2603 avdd.n234 avdd.n224 185
R2604 avdd.n233 avdd.n225 185
R2605 avdd.n28 avdd.n25 185
R2606 avdd.n243 avdd.n26 185
R2607 avdd.n211 avdd.n210 185
R2608 avdd.n212 avdd.n211 185
R2609 avdd.n39 avdd.n38 185
R2610 avdd.n206 avdd.n196 185
R2611 avdd.n205 avdd.n197 185
R2612 avdd.n36 avdd.n33 185
R2613 avdd.n215 avdd.n34 185
R2614 avdd.n183 avdd.n182 185
R2615 avdd.n184 avdd.n183 185
R2616 avdd.n47 avdd.n46 185
R2617 avdd.n178 avdd.n168 185
R2618 avdd.n177 avdd.n169 185
R2619 avdd.n44 avdd.n41 185
R2620 avdd.n187 avdd.n42 185
R2621 avdd.n155 avdd.n154 185
R2622 avdd.n156 avdd.n155 185
R2623 avdd.n55 avdd.n54 185
R2624 avdd.n150 avdd.n140 185
R2625 avdd.n149 avdd.n141 185
R2626 avdd.n52 avdd.n49 185
R2627 avdd.n159 avdd.n50 185
R2628 avdd.n127 avdd.n126 185
R2629 avdd.n128 avdd.n127 185
R2630 avdd.n63 avdd.n62 185
R2631 avdd.n122 avdd.n112 185
R2632 avdd.n121 avdd.n113 185
R2633 avdd.n60 avdd.n57 185
R2634 avdd.n131 avdd.n58 185
R2635 avdd.n76 avdd.n75 185
R2636 avdd.n71 avdd.n70 185
R2637 avdd.n70 avdd.n69 185
R2638 avdd.n92 avdd.n91 185
R2639 avdd.n93 avdd.n92 185
R2640 avdd.n72 avdd.n67 185
R2641 avdd.n94 avdd.n67 185
R2642 avdd.n96 avdd.n68 185
R2643 avdd.n96 avdd.n95 185
R2644 avdd.n97 avdd.n65 185
R2645 avdd.n98 avdd.n97 185
R2646 avdd.n103 avdd.n66 185
R2647 avdd.n99 avdd.n66 185
R2648 avdd.n102 avdd.n101 185
R2649 avdd.n101 avdd.n100 185
R2650 avdd.n659 avdd.n658 185
R2651 avdd.n660 avdd.n659 185
R2652 avdd.n343 avdd.n342 185
R2653 avdd.n654 avdd.n644 185
R2654 avdd.n653 avdd.n645 185
R2655 avdd.n340 avdd.n337 185
R2656 avdd.n663 avdd.n338 185
R2657 avdd.n631 avdd.n630 185
R2658 avdd.n632 avdd.n631 185
R2659 avdd.n351 avdd.n350 185
R2660 avdd.n626 avdd.n616 185
R2661 avdd.n625 avdd.n617 185
R2662 avdd.n348 avdd.n345 185
R2663 avdd.n635 avdd.n346 185
R2664 avdd.n603 avdd.n602 185
R2665 avdd.n604 avdd.n603 185
R2666 avdd.n359 avdd.n358 185
R2667 avdd.n598 avdd.n588 185
R2668 avdd.n597 avdd.n589 185
R2669 avdd.n356 avdd.n353 185
R2670 avdd.n607 avdd.n354 185
R2671 avdd.n575 avdd.n574 185
R2672 avdd.n576 avdd.n575 185
R2673 avdd.n367 avdd.n366 185
R2674 avdd.n570 avdd.n560 185
R2675 avdd.n569 avdd.n561 185
R2676 avdd.n364 avdd.n361 185
R2677 avdd.n579 avdd.n362 185
R2678 avdd.n547 avdd.n546 185
R2679 avdd.n548 avdd.n547 185
R2680 avdd.n375 avdd.n374 185
R2681 avdd.n542 avdd.n532 185
R2682 avdd.n541 avdd.n533 185
R2683 avdd.n372 avdd.n369 185
R2684 avdd.n551 avdd.n370 185
R2685 avdd.n519 avdd.n518 185
R2686 avdd.n520 avdd.n519 185
R2687 avdd.n383 avdd.n382 185
R2688 avdd.n514 avdd.n504 185
R2689 avdd.n513 avdd.n505 185
R2690 avdd.n380 avdd.n377 185
R2691 avdd.n523 avdd.n378 185
R2692 avdd.n491 avdd.n490 185
R2693 avdd.n492 avdd.n491 185
R2694 avdd.n391 avdd.n390 185
R2695 avdd.n486 avdd.n476 185
R2696 avdd.n485 avdd.n477 185
R2697 avdd.n388 avdd.n385 185
R2698 avdd.n495 avdd.n386 185
R2699 avdd.n463 avdd.n462 185
R2700 avdd.n464 avdd.n463 185
R2701 avdd.n399 avdd.n398 185
R2702 avdd.n458 avdd.n448 185
R2703 avdd.n457 avdd.n449 185
R2704 avdd.n396 avdd.n393 185
R2705 avdd.n467 avdd.n394 185
R2706 avdd.n412 avdd.n411 185
R2707 avdd.n407 avdd.n406 185
R2708 avdd.n406 avdd.n405 185
R2709 avdd.n428 avdd.n427 185
R2710 avdd.n429 avdd.n428 185
R2711 avdd.n408 avdd.n403 185
R2712 avdd.n430 avdd.n403 185
R2713 avdd.n432 avdd.n404 185
R2714 avdd.n432 avdd.n431 185
R2715 avdd.n433 avdd.n401 185
R2716 avdd.n434 avdd.n433 185
R2717 avdd.n439 avdd.n402 185
R2718 avdd.n435 avdd.n402 185
R2719 avdd.n438 avdd.n437 185
R2720 avdd.n437 avdd.n436 185
R2721 avdd.n679 avdd.n677 185
R2722 avdd.n680 avdd.n679 185
R2723 avdd.n683 avdd.n678 185
R2724 avdd.n924 avdd.n923 185
R2725 avdd.n923 avdd.n922 185
R2726 avdd.n703 avdd.n702 185
R2727 avdd.n921 avdd.n703 185
R2728 avdd.n919 avdd.n918 185
R2729 avdd.n920 avdd.n919 185
R2730 avdd.n913 avdd.n912 185
R2731 avdd.n912 avdd.n706 185
R2732 avdd.n911 avdd.n709 185
R2733 avdd.n911 avdd.n910 185
R2734 avdd.n712 avdd.n710 185
R2735 avdd.n909 avdd.n710 185
R2736 avdd.n907 avdd.n906 185
R2737 avdd.n908 avdd.n907 185
R2738 avdd.n905 avdd.n711 185
R2739 avdd.n723 avdd.n711 185
R2740 avdd.n724 avdd.n718 185
R2741 avdd.n725 avdd.n724 185
R2742 avdd.n899 avdd.n898 185
R2743 avdd.n898 avdd.n897 185
R2744 avdd.n722 avdd.n721 185
R2745 avdd.n896 avdd.n722 185
R2746 avdd.n894 avdd.n893 185
R2747 avdd.n895 avdd.n894 185
R2748 avdd.n888 avdd.n887 185
R2749 avdd.n887 avdd.n726 185
R2750 avdd.n886 avdd.n729 185
R2751 avdd.n886 avdd.n885 185
R2752 avdd.n732 avdd.n730 185
R2753 avdd.n884 avdd.n730 185
R2754 avdd.n882 avdd.n881 185
R2755 avdd.n883 avdd.n882 185
R2756 avdd.n880 avdd.n731 185
R2757 avdd.n743 avdd.n731 185
R2758 avdd.n744 avdd.n738 185
R2759 avdd.n745 avdd.n744 185
R2760 avdd.n874 avdd.n873 185
R2761 avdd.n873 avdd.n872 185
R2762 avdd.n742 avdd.n741 185
R2763 avdd.n871 avdd.n742 185
R2764 avdd.n869 avdd.n868 185
R2765 avdd.n870 avdd.n869 185
R2766 avdd.n863 avdd.n862 185
R2767 avdd.n862 avdd.n746 185
R2768 avdd.n861 avdd.n749 185
R2769 avdd.n861 avdd.n860 185
R2770 avdd.n752 avdd.n750 185
R2771 avdd.n859 avdd.n750 185
R2772 avdd.n857 avdd.n856 185
R2773 avdd.n858 avdd.n857 185
R2774 avdd.n855 avdd.n751 185
R2775 avdd.n763 avdd.n751 185
R2776 avdd.n764 avdd.n758 185
R2777 avdd.n765 avdd.n764 185
R2778 avdd.n849 avdd.n848 185
R2779 avdd.n848 avdd.n847 185
R2780 avdd.n762 avdd.n761 185
R2781 avdd.n846 avdd.n762 185
R2782 avdd.n844 avdd.n843 185
R2783 avdd.n845 avdd.n844 185
R2784 avdd.n838 avdd.n837 185
R2785 avdd.n837 avdd.n766 185
R2786 avdd.n836 avdd.n769 185
R2787 avdd.n836 avdd.n835 185
R2788 avdd.n772 avdd.n770 185
R2789 avdd.n834 avdd.n770 185
R2790 avdd.n832 avdd.n831 185
R2791 avdd.n833 avdd.n832 185
R2792 avdd.n830 avdd.n771 185
R2793 avdd.n783 avdd.n771 185
R2794 avdd.n784 avdd.n778 185
R2795 avdd.n785 avdd.n784 185
R2796 avdd.n824 avdd.n823 185
R2797 avdd.n823 avdd.n822 185
R2798 avdd.n782 avdd.n781 185
R2799 avdd.n821 avdd.n782 185
R2800 avdd.n819 avdd.n818 185
R2801 avdd.n820 avdd.n819 185
R2802 avdd.n813 avdd.n812 185
R2803 avdd.n812 avdd.n786 185
R2804 avdd.n811 avdd.n789 185
R2805 avdd.n811 avdd.n810 185
R2806 avdd.n792 avdd.n790 185
R2807 avdd.n809 avdd.n790 185
R2808 avdd.n807 avdd.n806 185
R2809 avdd.n808 avdd.n807 185
R2810 avdd.n805 avdd.n791 185
R2811 avdd.n931 avdd.n697 185
R2812 avdd.n930 avdd.n698 185
R2813 avdd.n704 avdd.n698 185
R2814 avdd.n929 avdd.n699 185
R2815 avdd.n705 avdd.n699 185
R2816 avdd.n1126 avdd.t246 180.231
R2817 avdd.n1166 avdd.t227 180.231
R2818 avdd.n1372 avdd.t240 180.231
R2819 avdd.n1412 avdd.t236 180.231
R2820 avdd.n705 avdd.n704 175.386
R2821 avdd.n921 avdd.n920 175.386
R2822 avdd.n910 avdd.n909 175.386
R2823 avdd.n725 avdd.n723 175.386
R2824 avdd.n896 avdd.n895 175.386
R2825 avdd.n885 avdd.n884 175.386
R2826 avdd.n745 avdd.n743 175.386
R2827 avdd.n871 avdd.n870 175.386
R2828 avdd.n860 avdd.n859 175.386
R2829 avdd.n765 avdd.n763 175.386
R2830 avdd.n846 avdd.n845 175.386
R2831 avdd.n835 avdd.n834 175.386
R2832 avdd.n785 avdd.n783 175.386
R2833 avdd.n821 avdd.n820 175.386
R2834 avdd.n810 avdd.n809 175.386
R2835 avdd.n922 avdd.t530 169.905
R2836 avdd.t46 avdd.n706 169.905
R2837 avdd.n908 avdd.t408 169.905
R2838 avdd.n897 avdd.t104 169.905
R2839 avdd.t157 avdd.n726 169.905
R2840 avdd.n883 avdd.t577 169.905
R2841 avdd.n872 avdd.t539 169.905
R2842 avdd.t609 avdd.n746 169.905
R2843 avdd.n858 avdd.t207 169.905
R2844 avdd.n847 avdd.t118 169.905
R2845 avdd.t579 avdd.n766 169.905
R2846 avdd.n833 avdd.t581 169.905
R2847 avdd.n822 avdd.t106 169.905
R2848 avdd.t211 avdd.n786 169.905
R2849 avdd.n808 avdd.t532 169.905
R2850 avdd.t574 avdd.n1535 167.023
R2851 avdd.n1589 avdd.n1588 165.936
R2852 avdd.n1591 avdd.n1590 155.859
R2853 avdd.n1595 avdd.n1594 155.859
R2854 avdd.n1160 avdd.t22 155.153
R2855 avdd.n1160 avdd.t18 155.153
R2856 avdd.n1406 avdd.t133 155.153
R2857 avdd.n1406 avdd.t125 155.153
R2858 avdd.t324 avdd.t574 153.764
R2859 avdd.n312 avdd.n311 153.571
R2860 avdd.n284 avdd.n283 153.571
R2861 avdd.n256 avdd.n255 153.571
R2862 avdd.n228 avdd.n227 153.571
R2863 avdd.n200 avdd.n199 153.571
R2864 avdd.n172 avdd.n171 153.571
R2865 avdd.n144 avdd.n143 153.571
R2866 avdd.n116 avdd.n115 153.571
R2867 avdd.n83 avdd.n82 153.571
R2868 avdd.n648 avdd.n647 153.571
R2869 avdd.n620 avdd.n619 153.571
R2870 avdd.n592 avdd.n591 153.571
R2871 avdd.n564 avdd.n563 153.571
R2872 avdd.n536 avdd.n535 153.571
R2873 avdd.n508 avdd.n507 153.571
R2874 avdd.n480 avdd.n479 153.571
R2875 avdd.n452 avdd.n451 153.571
R2876 avdd.n419 avdd.n418 153.571
R2877 avdd.t58 avdd.n1631 149.893
R2878 avdd.n1633 avdd.t78 149.893
R2879 avdd.t492 avdd.n1646 149.893
R2880 avdd.n1647 avdd.t413 149.893
R2881 avdd.n1634 avdd.n1628 125.742
R2882 avdd.n1626 avdd.n1609 125.742
R2883 avdd.t557 avdd.t218 121.877
R2884 avdd.t545 avdd.t555 121.877
R2885 avdd.n93 avdd.n69 120.317
R2886 avdd.n95 avdd.n94 120.317
R2887 avdd.n99 avdd.n98 120.317
R2888 avdd.n100 avdd.n99 120.317
R2889 avdd.n431 avdd.n430 120.317
R2890 avdd.n435 avdd.n434 120.317
R2891 avdd.n436 avdd.n435 120.317
R2892 avdd.n429 avdd.n405 119.064
R2893 avdd.n1122 avdd.t426 116.782
R2894 avdd.n1122 avdd.t436 116.782
R2895 avdd.n1368 avdd.t590 116.782
R2896 avdd.n1368 avdd.t598 116.782
R2897 avdd.t72 avdd.t58 110.959
R2898 avdd.t88 avdd.t72 110.959
R2899 avdd.t68 avdd.t88 110.959
R2900 avdd.t84 avdd.t68 110.959
R2901 avdd.t80 avdd.t84 110.959
R2902 avdd.t62 avdd.t80 110.959
R2903 avdd.t76 avdd.t62 110.959
R2904 avdd.t74 avdd.t60 110.959
R2905 avdd.t70 avdd.t74 110.959
R2906 avdd.t86 avdd.t70 110.959
R2907 avdd.t66 avdd.t86 110.959
R2908 avdd.t82 avdd.t66 110.959
R2909 avdd.t64 avdd.t82 110.959
R2910 avdd.t78 avdd.t64 110.959
R2911 avdd.t491 avdd.t492 110.959
R2912 avdd.t310 avdd.t491 110.959
R2913 avdd.t156 avdd.t310 110.959
R2914 avdd.t155 avdd.t156 110.959
R2915 avdd.t249 avdd.t155 110.959
R2916 avdd.t180 avdd.t249 110.959
R2917 avdd.t179 avdd.t180 110.959
R2918 avdd.t339 avdd.t179 110.959
R2919 avdd.t504 avdd.t339 110.959
R2920 avdd.t503 avdd.t504 110.959
R2921 avdd.t281 avdd.t503 110.959
R2922 avdd.t522 avdd.t281 110.959
R2923 avdd.t523 avdd.t522 110.959
R2924 avdd.t381 avdd.t523 110.959
R2925 avdd.t109 avdd.t381 110.959
R2926 avdd.t108 avdd.t109 110.959
R2927 avdd.t268 avdd.t108 110.959
R2928 avdd.t152 avdd.t268 110.959
R2929 avdd.t151 avdd.t152 110.959
R2930 avdd.t399 avdd.t151 110.959
R2931 avdd.t420 avdd.t399 110.959
R2932 avdd.t419 avdd.t420 110.959
R2933 avdd.t387 avdd.t419 110.959
R2934 avdd.t170 avdd.t387 110.959
R2935 avdd.t171 avdd.t170 110.959
R2936 avdd.t374 avdd.t171 110.959
R2937 avdd.t490 avdd.t374 110.959
R2938 avdd.t489 avdd.t490 110.959
R2939 avdd.t385 avdd.t489 110.959
R2940 avdd.t167 avdd.t385 110.959
R2941 avdd.t168 avdd.t167 110.959
R2942 avdd.t303 avdd.t168 110.959
R2943 avdd.t402 avdd.t303 110.959
R2944 avdd.t403 avdd.t402 110.959
R2945 avdd.t397 avdd.t403 110.959
R2946 avdd.t499 avdd.t397 110.959
R2947 avdd.t500 avdd.t499 110.959
R2948 avdd.t401 avdd.t500 110.959
R2949 avdd.t2 avdd.t401 110.959
R2950 avdd.t3 avdd.t2 110.959
R2951 avdd.t363 avdd.t3 110.959
R2952 avdd.t214 avdd.t363 110.959
R2953 avdd.t213 avdd.t214 110.959
R2954 avdd.t254 avdd.t213 110.959
R2955 avdd.t412 avdd.t254 110.959
R2956 avdd.t413 avdd.t412 110.959
R2957 avdd.n324 avdd.t159 106.817
R2958 avdd.n296 avdd.t519 106.817
R2959 avdd.n268 avdd.t452 106.817
R2960 avdd.n240 avdd.t584 106.817
R2961 avdd.n212 avdd.t404 106.817
R2962 avdd.n184 avdd.t120 106.817
R2963 avdd.n156 avdd.t513 106.817
R2964 avdd.n128 avdd.t486 106.817
R2965 avdd.n660 avdd.t416 106.817
R2966 avdd.n632 avdd.t496 106.817
R2967 avdd.n604 avdd.t440 106.817
R2968 avdd.n576 avdd.t535 106.817
R2969 avdd.n548 avdd.t114 106.817
R2970 avdd.n520 avdd.t56 106.817
R2971 avdd.n492 avdd.t607 106.817
R2972 avdd.n464 avdd.t12 106.817
R2973 avdd.t565 avdd.n93 106.531
R2974 avdd.t221 avdd.n429 106.531
R2975 avdd.n1163 avdd.n975 105.412
R2976 avdd.n1409 avdd.n1221 105.412
R2977 avdd.t159 avdd.t153 102.091
R2978 avdd.t519 avdd.t517 102.091
R2979 avdd.t452 avdd.t454 102.091
R2980 avdd.t584 avdd.t172 102.091
R2981 avdd.t404 avdd.t406 102.091
R2982 avdd.t120 avdd.t0 102.091
R2983 avdd.t513 avdd.t515 102.091
R2984 avdd.t486 avdd.t450 102.091
R2985 avdd.t416 avdd.t215 102.091
R2986 avdd.t496 avdd.t110 102.091
R2987 avdd.t440 avdd.t442 102.091
R2988 avdd.t535 avdd.t116 102.091
R2989 avdd.t114 avdd.t112 102.091
R2990 avdd.t56 avdd.t54 102.091
R2991 avdd.t607 avdd.t528 102.091
R2992 avdd.t12 avdd.t10 102.091
R2993 avdd.t165 avdd.n69 101.564
R2994 avdd.t48 avdd.n405 101.564
R2995 avdd.n969 avdd.n968 99.0123
R2996 avdd.n974 avdd.n973 99.0123
R2997 avdd.n1215 avdd.n1214 99.0123
R2998 avdd.n1220 avdd.n1219 99.0123
R2999 avdd.n100 avdd.t421 97.7578
R3000 avdd.n436 avdd.t102 97.7578
R3001 avdd.t569 avdd.n1517 96.5971
R3002 avdd.n1169 avdd.n1168 94.1181
R3003 avdd.n1129 avdd.n1128 94.1181
R3004 avdd.n1415 avdd.n1414 94.1181
R3005 avdd.n1375 avdd.n1374 94.1181
R3006 avdd.n1018 avdd.n1013 91.1064
R3007 avdd.n1264 avdd.n1259 91.1064
R3008 avdd.t96 avdd.t569 88.8801
R3009 avdd.n6 avdd.n3 86.068
R3010 avdd.n309 avdd.n5 86.068
R3011 avdd.n325 avdd.n2 86.068
R3012 avdd.n308 avdd.n3 86.068
R3013 avdd.n5 avdd.n4 86.068
R3014 avdd.n14 avdd.n11 86.068
R3015 avdd.n281 avdd.n13 86.068
R3016 avdd.n297 avdd.n10 86.068
R3017 avdd.n280 avdd.n11 86.068
R3018 avdd.n13 avdd.n12 86.068
R3019 avdd.n22 avdd.n19 86.068
R3020 avdd.n253 avdd.n21 86.068
R3021 avdd.n269 avdd.n18 86.068
R3022 avdd.n252 avdd.n19 86.068
R3023 avdd.n21 avdd.n20 86.068
R3024 avdd.n30 avdd.n27 86.068
R3025 avdd.n225 avdd.n29 86.068
R3026 avdd.n241 avdd.n26 86.068
R3027 avdd.n224 avdd.n27 86.068
R3028 avdd.n29 avdd.n28 86.068
R3029 avdd.n38 avdd.n35 86.068
R3030 avdd.n197 avdd.n37 86.068
R3031 avdd.n213 avdd.n34 86.068
R3032 avdd.n196 avdd.n35 86.068
R3033 avdd.n37 avdd.n36 86.068
R3034 avdd.n46 avdd.n43 86.068
R3035 avdd.n169 avdd.n45 86.068
R3036 avdd.n185 avdd.n42 86.068
R3037 avdd.n168 avdd.n43 86.068
R3038 avdd.n45 avdd.n44 86.068
R3039 avdd.n54 avdd.n51 86.068
R3040 avdd.n141 avdd.n53 86.068
R3041 avdd.n157 avdd.n50 86.068
R3042 avdd.n140 avdd.n51 86.068
R3043 avdd.n53 avdd.n52 86.068
R3044 avdd.n62 avdd.n59 86.068
R3045 avdd.n113 avdd.n61 86.068
R3046 avdd.n129 avdd.n58 86.068
R3047 avdd.n112 avdd.n59 86.068
R3048 avdd.n61 avdd.n60 86.068
R3049 avdd.n342 avdd.n339 86.068
R3050 avdd.n645 avdd.n341 86.068
R3051 avdd.n661 avdd.n338 86.068
R3052 avdd.n644 avdd.n339 86.068
R3053 avdd.n341 avdd.n340 86.068
R3054 avdd.n350 avdd.n347 86.068
R3055 avdd.n617 avdd.n349 86.068
R3056 avdd.n633 avdd.n346 86.068
R3057 avdd.n616 avdd.n347 86.068
R3058 avdd.n349 avdd.n348 86.068
R3059 avdd.n358 avdd.n355 86.068
R3060 avdd.n589 avdd.n357 86.068
R3061 avdd.n605 avdd.n354 86.068
R3062 avdd.n588 avdd.n355 86.068
R3063 avdd.n357 avdd.n356 86.068
R3064 avdd.n366 avdd.n363 86.068
R3065 avdd.n561 avdd.n365 86.068
R3066 avdd.n577 avdd.n362 86.068
R3067 avdd.n560 avdd.n363 86.068
R3068 avdd.n365 avdd.n364 86.068
R3069 avdd.n374 avdd.n371 86.068
R3070 avdd.n533 avdd.n373 86.068
R3071 avdd.n549 avdd.n370 86.068
R3072 avdd.n532 avdd.n371 86.068
R3073 avdd.n373 avdd.n372 86.068
R3074 avdd.n382 avdd.n379 86.068
R3075 avdd.n505 avdd.n381 86.068
R3076 avdd.n521 avdd.n378 86.068
R3077 avdd.n504 avdd.n379 86.068
R3078 avdd.n381 avdd.n380 86.068
R3079 avdd.n390 avdd.n387 86.068
R3080 avdd.n477 avdd.n389 86.068
R3081 avdd.n493 avdd.n386 86.068
R3082 avdd.n476 avdd.n387 86.068
R3083 avdd.n389 avdd.n388 86.068
R3084 avdd.n398 avdd.n395 86.068
R3085 avdd.n449 avdd.n397 86.068
R3086 avdd.n465 avdd.n394 86.068
R3087 avdd.n448 avdd.n395 86.068
R3088 avdd.n397 avdd.n396 86.068
R3089 avdd.n681 avdd.n678 86.068
R3090 avdd.n798 avdd.t532 82.3568
R3091 avdd.t545 avdd.t100 73.4459
R3092 avdd.n95 avdd.t52 72.6918
R3093 avdd.n431 avdd.t8 72.6918
R3094 avdd.n968 avdd.n956 71.5299
R3095 avdd.n975 avdd.n974 71.5299
R3096 avdd.n1214 avdd.n1202 71.5299
R3097 avdd.n1221 avdd.n1220 71.5299
R3098 avdd.t547 avdd.n1538 69.9865
R3099 avdd.n798 avdd.n791 68.6629
R3100 avdd.n1544 avdd.t164 59.3422
R3101 avdd.t231 avdd.t557 58.0117
R3102 avdd.n1632 avdd.t76 55.4795
R3103 avdd.t60 avdd.n1632 55.4795
R3104 avdd.n1624 avdd.t79 54.6604
R3105 avdd.n1607 avdd.t59 54.6604
R3106 avdd.n1527 avdd.t570 53.8832
R3107 avdd.n1521 avdd.t548 53.8832
R3108 avdd.n1520 avdd.t575 53.8832
R3109 avdd.n1505 avdd.n1504 50.4475
R3110 avdd.n1567 avdd.t335 49.5908
R3111 avdd.n1551 avdd.t335 49.5908
R3112 avdd.n324 avdd.n3 49.4675
R3113 avdd.n324 avdd.n5 49.4675
R3114 avdd.n325 avdd.n324 49.4675
R3115 avdd.n296 avdd.n11 49.4675
R3116 avdd.n296 avdd.n13 49.4675
R3117 avdd.n297 avdd.n296 49.4675
R3118 avdd.n268 avdd.n19 49.4675
R3119 avdd.n268 avdd.n21 49.4675
R3120 avdd.n269 avdd.n268 49.4675
R3121 avdd.n240 avdd.n27 49.4675
R3122 avdd.n240 avdd.n29 49.4675
R3123 avdd.n241 avdd.n240 49.4675
R3124 avdd.n212 avdd.n35 49.4675
R3125 avdd.n212 avdd.n37 49.4675
R3126 avdd.n213 avdd.n212 49.4675
R3127 avdd.n184 avdd.n43 49.4675
R3128 avdd.n184 avdd.n45 49.4675
R3129 avdd.n185 avdd.n184 49.4675
R3130 avdd.n156 avdd.n51 49.4675
R3131 avdd.n156 avdd.n53 49.4675
R3132 avdd.n157 avdd.n156 49.4675
R3133 avdd.n128 avdd.n59 49.4675
R3134 avdd.n128 avdd.n61 49.4675
R3135 avdd.n129 avdd.n128 49.4675
R3136 avdd.n660 avdd.n339 49.4675
R3137 avdd.n660 avdd.n341 49.4675
R3138 avdd.n661 avdd.n660 49.4675
R3139 avdd.n632 avdd.n347 49.4675
R3140 avdd.n632 avdd.n349 49.4675
R3141 avdd.n633 avdd.n632 49.4675
R3142 avdd.n604 avdd.n355 49.4675
R3143 avdd.n604 avdd.n357 49.4675
R3144 avdd.n605 avdd.n604 49.4675
R3145 avdd.n576 avdd.n363 49.4675
R3146 avdd.n576 avdd.n365 49.4675
R3147 avdd.n577 avdd.n576 49.4675
R3148 avdd.n548 avdd.n371 49.4675
R3149 avdd.n548 avdd.n373 49.4675
R3150 avdd.n549 avdd.n548 49.4675
R3151 avdd.n520 avdd.n379 49.4675
R3152 avdd.n520 avdd.n381 49.4675
R3153 avdd.n521 avdd.n520 49.4675
R3154 avdd.n492 avdd.n387 49.4675
R3155 avdd.n492 avdd.n389 49.4675
R3156 avdd.n493 avdd.n492 49.4675
R3157 avdd.n464 avdd.n395 49.4675
R3158 avdd.n464 avdd.n397 49.4675
R3159 avdd.n465 avdd.n464 49.4675
R3160 avdd.n681 avdd.n680 49.4675
R3161 avdd.n1623 avdd.n1622 49.1214
R3162 avdd.n1621 avdd.n1620 49.1214
R3163 avdd.n1619 avdd.n1618 49.1214
R3164 avdd.n1617 avdd.n1616 49.1214
R3165 avdd.n1615 avdd.n1614 49.1214
R3166 avdd.n1613 avdd.n1612 49.1214
R3167 avdd.n1611 avdd.n1610 49.1214
R3168 avdd.t218 avdd.t100 48.4319
R3169 avdd.n1529 avdd.n1528 48.3442
R3170 avdd.n1531 avdd.n1530 48.3442
R3171 avdd.n1556 avdd.n1555 48.2034
R3172 avdd.n1558 avdd.n1557 48.2034
R3173 avdd.n1564 avdd.n1563 48.2034
R3174 avdd.n1571 avdd.n1570 48.2034
R3175 avdd.n1573 avdd.n1572 48.2034
R3176 avdd.n1575 avdd.n1574 48.2034
R3177 avdd.n1577 avdd.n1576 48.2034
R3178 avdd.n1553 avdd.t266 48.0365
R3179 avdd.n1578 avdd.t232 48.0365
R3180 avdd.n98 avdd.t52 47.6258
R3181 avdd.n434 avdd.t8 47.6258
R3182 avdd.t163 avdd.t220 47.3674
R3183 avdd.t220 avdd.t234 47.3674
R3184 avdd.t234 avdd.t217 47.3674
R3185 avdd.t351 avdd.t217 47.3674
R3186 avdd.t344 avdd.t573 47.3674
R3187 avdd.t571 avdd.t344 47.3674
R3188 avdd.t164 avdd.t571 47.3674
R3189 avdd.n1170 avdd.n1169 44.8005
R3190 avdd.n1130 avdd.n1129 44.8005
R3191 avdd.n1416 avdd.n1415 44.8005
R3192 avdd.n1376 avdd.n1375 44.8005
R3193 avdd.n1019 avdd.n1014 43.2946
R3194 avdd.n1265 avdd.n1260 43.2946
R3195 avdd.n1517 avdd.t446 42.8436
R3196 avdd.n1560 avdd.n1559 42.4975
R3197 avdd.n1562 avdd.n1552 42.4505
R3198 avdd.n1584 avdd.t547 41.247
R3199 avdd.n1538 avdd.t231 38.5859
R3200 avdd.n973 avdd.n972 37.0005
R3201 avdd.n970 avdd.n969 37.0005
R3202 avdd.n1219 avdd.n1218 37.0005
R3203 avdd.n1216 avdd.n1215 37.0005
R3204 avdd.n1483 avdd.n1482 36.4934
R3205 avdd.n322 avdd.n7 36.1417
R3206 avdd.n318 avdd.n7 36.1417
R3207 avdd.n318 avdd.n317 36.1417
R3208 avdd.n317 avdd.n1 36.1417
R3209 avdd.n327 avdd.n1 36.1417
R3210 avdd.n327 avdd.n326 36.1417
R3211 avdd.n294 avdd.n15 36.1417
R3212 avdd.n290 avdd.n15 36.1417
R3213 avdd.n290 avdd.n289 36.1417
R3214 avdd.n289 avdd.n9 36.1417
R3215 avdd.n299 avdd.n9 36.1417
R3216 avdd.n299 avdd.n298 36.1417
R3217 avdd.n266 avdd.n23 36.1417
R3218 avdd.n262 avdd.n23 36.1417
R3219 avdd.n262 avdd.n261 36.1417
R3220 avdd.n261 avdd.n17 36.1417
R3221 avdd.n271 avdd.n17 36.1417
R3222 avdd.n271 avdd.n270 36.1417
R3223 avdd.n238 avdd.n31 36.1417
R3224 avdd.n234 avdd.n31 36.1417
R3225 avdd.n234 avdd.n233 36.1417
R3226 avdd.n233 avdd.n25 36.1417
R3227 avdd.n243 avdd.n25 36.1417
R3228 avdd.n243 avdd.n242 36.1417
R3229 avdd.n210 avdd.n39 36.1417
R3230 avdd.n206 avdd.n39 36.1417
R3231 avdd.n206 avdd.n205 36.1417
R3232 avdd.n205 avdd.n33 36.1417
R3233 avdd.n215 avdd.n33 36.1417
R3234 avdd.n215 avdd.n214 36.1417
R3235 avdd.n182 avdd.n47 36.1417
R3236 avdd.n178 avdd.n47 36.1417
R3237 avdd.n178 avdd.n177 36.1417
R3238 avdd.n177 avdd.n41 36.1417
R3239 avdd.n187 avdd.n41 36.1417
R3240 avdd.n187 avdd.n186 36.1417
R3241 avdd.n154 avdd.n55 36.1417
R3242 avdd.n150 avdd.n55 36.1417
R3243 avdd.n150 avdd.n149 36.1417
R3244 avdd.n149 avdd.n49 36.1417
R3245 avdd.n159 avdd.n49 36.1417
R3246 avdd.n159 avdd.n158 36.1417
R3247 avdd.n126 avdd.n63 36.1417
R3248 avdd.n122 avdd.n63 36.1417
R3249 avdd.n122 avdd.n121 36.1417
R3250 avdd.n121 avdd.n57 36.1417
R3251 avdd.n131 avdd.n57 36.1417
R3252 avdd.n131 avdd.n130 36.1417
R3253 avdd.n76 avdd.n71 36.1417
R3254 avdd.n91 avdd.n71 36.1417
R3255 avdd.n91 avdd.n72 36.1417
R3256 avdd.n72 avdd.n68 36.1417
R3257 avdd.n68 avdd.n65 36.1417
R3258 avdd.n103 avdd.n65 36.1417
R3259 avdd.n103 avdd.n102 36.1417
R3260 avdd.n658 avdd.n343 36.1417
R3261 avdd.n654 avdd.n343 36.1417
R3262 avdd.n654 avdd.n653 36.1417
R3263 avdd.n653 avdd.n337 36.1417
R3264 avdd.n663 avdd.n337 36.1417
R3265 avdd.n663 avdd.n662 36.1417
R3266 avdd.n630 avdd.n351 36.1417
R3267 avdd.n626 avdd.n351 36.1417
R3268 avdd.n626 avdd.n625 36.1417
R3269 avdd.n625 avdd.n345 36.1417
R3270 avdd.n635 avdd.n345 36.1417
R3271 avdd.n635 avdd.n634 36.1417
R3272 avdd.n602 avdd.n359 36.1417
R3273 avdd.n598 avdd.n359 36.1417
R3274 avdd.n598 avdd.n597 36.1417
R3275 avdd.n597 avdd.n353 36.1417
R3276 avdd.n607 avdd.n353 36.1417
R3277 avdd.n607 avdd.n606 36.1417
R3278 avdd.n574 avdd.n367 36.1417
R3279 avdd.n570 avdd.n367 36.1417
R3280 avdd.n570 avdd.n569 36.1417
R3281 avdd.n569 avdd.n361 36.1417
R3282 avdd.n579 avdd.n361 36.1417
R3283 avdd.n579 avdd.n578 36.1417
R3284 avdd.n546 avdd.n375 36.1417
R3285 avdd.n542 avdd.n375 36.1417
R3286 avdd.n542 avdd.n541 36.1417
R3287 avdd.n541 avdd.n369 36.1417
R3288 avdd.n551 avdd.n369 36.1417
R3289 avdd.n551 avdd.n550 36.1417
R3290 avdd.n518 avdd.n383 36.1417
R3291 avdd.n514 avdd.n383 36.1417
R3292 avdd.n514 avdd.n513 36.1417
R3293 avdd.n513 avdd.n377 36.1417
R3294 avdd.n523 avdd.n377 36.1417
R3295 avdd.n523 avdd.n522 36.1417
R3296 avdd.n490 avdd.n391 36.1417
R3297 avdd.n486 avdd.n391 36.1417
R3298 avdd.n486 avdd.n485 36.1417
R3299 avdd.n485 avdd.n385 36.1417
R3300 avdd.n495 avdd.n385 36.1417
R3301 avdd.n495 avdd.n494 36.1417
R3302 avdd.n462 avdd.n399 36.1417
R3303 avdd.n458 avdd.n399 36.1417
R3304 avdd.n458 avdd.n457 36.1417
R3305 avdd.n457 avdd.n393 36.1417
R3306 avdd.n467 avdd.n393 36.1417
R3307 avdd.n467 avdd.n466 36.1417
R3308 avdd.n412 avdd.n407 36.1417
R3309 avdd.n427 avdd.n408 36.1417
R3310 avdd.n408 avdd.n404 36.1417
R3311 avdd.n404 avdd.n401 36.1417
R3312 avdd.n439 avdd.n401 36.1417
R3313 avdd.n439 avdd.n438 36.1417
R3314 avdd.n683 avdd.n677 36.1417
R3315 avdd.n683 avdd.n682 36.1417
R3316 avdd.n806 avdd.n805 36.1417
R3317 avdd.n805 avdd.n799 36.1417
R3318 avdd.n813 avdd.n789 36.1417
R3319 avdd.n792 avdd.n789 36.1417
R3320 avdd.n824 avdd.n781 36.1417
R3321 avdd.n818 avdd.n781 36.1417
R3322 avdd.n831 avdd.n830 36.1417
R3323 avdd.n830 avdd.n778 36.1417
R3324 avdd.n838 avdd.n769 36.1417
R3325 avdd.n772 avdd.n769 36.1417
R3326 avdd.n849 avdd.n761 36.1417
R3327 avdd.n843 avdd.n761 36.1417
R3328 avdd.n856 avdd.n855 36.1417
R3329 avdd.n855 avdd.n758 36.1417
R3330 avdd.n863 avdd.n749 36.1417
R3331 avdd.n752 avdd.n749 36.1417
R3332 avdd.n874 avdd.n741 36.1417
R3333 avdd.n868 avdd.n741 36.1417
R3334 avdd.n881 avdd.n880 36.1417
R3335 avdd.n880 avdd.n738 36.1417
R3336 avdd.n888 avdd.n729 36.1417
R3337 avdd.n732 avdd.n729 36.1417
R3338 avdd.n899 avdd.n721 36.1417
R3339 avdd.n893 avdd.n721 36.1417
R3340 avdd.n906 avdd.n905 36.1417
R3341 avdd.n905 avdd.n718 36.1417
R3342 avdd.n913 avdd.n709 36.1417
R3343 avdd.n712 avdd.n709 36.1417
R3344 avdd.n924 avdd.n702 36.1417
R3345 avdd.n918 avdd.n702 36.1417
R3346 avdd.n931 avdd.n930 36.1417
R3347 avdd.n930 avdd.n929 36.1417
R3348 avdd.n427 avdd.n407 35.7652
R3349 avdd.t555 avdd.t96 32.9977
R3350 avdd.n1525 avdd.n1513 31.624
R3351 avdd.n1536 avdd.n1533 31.624
R3352 avdd.n1601 avdd.n1508 31.624
R3353 avdd.n1119 avdd.n1041 31.2476
R3354 avdd.n1039 avdd.n1038 31.2476
R3355 avdd.n1365 avdd.n1287 31.2476
R3356 avdd.n1285 avdd.n1284 31.2476
R3357 avdd.n1482 avdd.n1455 31.2285
R3358 avdd.n1128 avdd.n1127 30.8338
R3359 avdd.n1127 avdd.n1126 30.8338
R3360 avdd.n1168 avdd.n1167 30.8338
R3361 avdd.n1167 avdd.n1166 30.8338
R3362 avdd.n1041 avdd.n1037 30.8338
R3363 avdd.n1039 avdd.n1036 30.8338
R3364 avdd.n1374 avdd.n1373 30.8338
R3365 avdd.n1373 avdd.n1372 30.8338
R3366 avdd.n1414 avdd.n1413 30.8338
R3367 avdd.n1413 avdd.n1412 30.8338
R3368 avdd.n1287 avdd.n1283 30.8338
R3369 avdd.n1285 avdd.n1282 30.8338
R3370 avdd.n1464 avdd.n1462 30.3029
R3371 avdd.n1488 avdd.n1483 27.9872
R3372 avdd.n1060 avdd.t187 27.6955
R3373 avdd.n1060 avdd.t19 27.6955
R3374 avdd.n1058 avdd.t190 27.6955
R3375 avdd.n1058 avdd.t21 27.6955
R3376 avdd.n1056 avdd.t188 27.6955
R3377 avdd.n1056 avdd.t20 27.6955
R3378 avdd.n1054 avdd.t196 27.6955
R3379 avdd.n1054 avdd.t32 27.6955
R3380 avdd.n1052 avdd.t40 27.6955
R3381 avdd.n1052 avdd.t191 27.6955
R3382 avdd.n1050 avdd.t41 27.6955
R3383 avdd.n1050 avdd.t192 27.6955
R3384 avdd.n1048 avdd.t44 27.6955
R3385 avdd.n1048 avdd.t194 27.6955
R3386 avdd.n1046 avdd.t42 27.6955
R3387 avdd.n1046 avdd.t193 27.6955
R3388 avdd.n1044 avdd.t23 27.6955
R3389 avdd.n1044 avdd.t197 27.6955
R3390 avdd.n1042 avdd.t45 27.6955
R3391 avdd.n1042 avdd.t195 27.6955
R3392 avdd.n981 avdd.t24 27.6955
R3393 avdd.n981 avdd.t199 27.6955
R3394 avdd.n1155 avdd.t30 27.6955
R3395 avdd.n1155 avdd.t182 27.6955
R3396 avdd.t283 avdd.n1104 27.6955
R3397 avdd.n1104 avdd.t198 27.6955
R3398 avdd.n1101 avdd.t290 27.6955
R3399 avdd.n1101 avdd.t201 27.6955
R3400 avdd.n1098 avdd.t288 27.6955
R3401 avdd.n1098 avdd.t200 27.6955
R3402 avdd.t353 avdd.n1093 27.6955
R3403 avdd.n1093 avdd.t184 27.6955
R3404 avdd.t367 avdd.n1090 27.6955
R3405 avdd.n1090 avdd.t26 27.6955
R3406 avdd.n1087 avdd.t369 27.6955
R3407 avdd.n1087 avdd.t27 27.6955
R3408 avdd.n1084 avdd.t383 27.6955
R3409 avdd.n1084 avdd.t29 27.6955
R3410 avdd.t376 avdd.n1079 27.6955
R3411 avdd.n1079 avdd.t28 27.6955
R3412 avdd.t247 avdd.n1076 27.6955
R3413 avdd.n1076 avdd.t36 27.6955
R3414 avdd.n1073 avdd.t392 27.6955
R3415 avdd.n1073 avdd.t31 27.6955
R3416 avdd.n1070 avdd.t256 27.6955
R3417 avdd.n1070 avdd.t38 27.6955
R3418 avdd.n1134 avdd.t274 27.6955
R3419 avdd.n1134 avdd.t39 27.6955
R3420 avdd.n986 avdd.t34 27.6955
R3421 avdd.n986 avdd.t251 27.6955
R3422 avdd.n988 avdd.t37 27.6955
R3423 avdd.n988 avdd.t261 27.6955
R3424 avdd.n990 avdd.t35 27.6955
R3425 avdd.n990 avdd.t258 27.6955
R3426 avdd.n992 avdd.t43 27.6955
R3427 avdd.n992 avdd.t295 27.6955
R3428 avdd.n994 avdd.t202 27.6955
R3429 avdd.n994 avdd.t315 27.6955
R3430 avdd.n996 avdd.t203 27.6955
R3431 avdd.n996 avdd.t318 27.6955
R3432 avdd.n998 avdd.t181 27.6955
R3433 avdd.n998 avdd.t333 27.6955
R3434 avdd.n1000 avdd.t204 27.6955
R3435 avdd.n1000 avdd.t328 27.6955
R3436 avdd.n1002 avdd.t185 27.6955
R3437 avdd.n1002 avdd.t389 27.6955
R3438 avdd.n1004 avdd.t183 27.6955
R3439 avdd.n1004 avdd.t341 27.6955
R3440 avdd.n1006 avdd.t186 27.6955
R3441 avdd.n1006 avdd.t394 27.6955
R3442 avdd.n1009 avdd.t189 27.6955
R3443 avdd.n1009 avdd.t228 27.6955
R3444 avdd.n1110 avdd.t425 27.6955
R3445 avdd.n1110 avdd.t435 27.6955
R3446 avdd.n1112 avdd.t433 27.6955
R3447 avdd.n1112 avdd.t427 27.6955
R3448 avdd.n1114 avdd.t437 27.6955
R3449 avdd.n1114 avdd.t429 27.6955
R3450 avdd.n1116 avdd.t439 27.6955
R3451 avdd.n1116 avdd.t178 27.6955
R3452 avdd.n1306 avdd.t137 27.6955
R3453 avdd.n1306 avdd.t480 27.6955
R3454 avdd.n1304 avdd.t135 27.6955
R3455 avdd.n1304 avdd.t478 27.6955
R3456 avdd.n1302 avdd.t136 27.6955
R3457 avdd.n1302 avdd.t479 27.6955
R3458 avdd.n1300 avdd.t134 27.6955
R3459 avdd.n1300 avdd.t477 27.6955
R3460 avdd.n1298 avdd.t462 27.6955
R3461 avdd.n1298 avdd.t131 27.6955
R3462 avdd.n1296 avdd.t472 27.6955
R3463 avdd.n1296 avdd.t139 27.6955
R3464 avdd.n1294 avdd.t460 27.6955
R3465 avdd.n1294 avdd.t130 27.6955
R3466 avdd.n1292 avdd.t471 27.6955
R3467 avdd.n1292 avdd.t129 27.6955
R3468 avdd.n1290 avdd.t470 27.6955
R3469 avdd.n1290 avdd.t128 27.6955
R3470 avdd.n1288 avdd.t469 27.6955
R3471 avdd.n1288 avdd.t126 27.6955
R3472 avdd.n1227 avdd.t459 27.6955
R3473 avdd.n1227 avdd.t148 27.6955
R3474 avdd.n1401 avdd.t481 27.6955
R3475 avdd.n1401 avdd.t142 27.6955
R3476 avdd.t365 avdd.n1350 27.6955
R3477 avdd.n1350 avdd.t145 27.6955
R3478 avdd.n1347 avdd.t349 27.6955
R3479 avdd.n1347 avdd.t143 27.6955
R3480 avdd.n1344 avdd.t355 27.6955
R3481 avdd.n1344 avdd.t144 27.6955
R3482 avdd.t347 avdd.n1339 27.6955
R3483 avdd.n1339 avdd.t141 27.6955
R3484 avdd.t276 avdd.n1336 27.6955
R3485 avdd.n1336 avdd.t468 27.6955
R3486 avdd.n1333 avdd.t331 27.6955
R3487 avdd.n1333 avdd.t476 27.6955
R3488 avdd.n1330 avdd.t272 27.6955
R3489 avdd.n1330 avdd.t467 27.6955
R3490 avdd.t326 avdd.n1325 27.6955
R3491 avdd.n1325 avdd.t475 27.6955
R3492 avdd.t308 avdd.n1322 27.6955
R3493 avdd.n1322 avdd.t474 27.6955
R3494 avdd.n1319 avdd.t301 27.6955
R3495 avdd.n1319 avdd.t473 27.6955
R3496 avdd.n1316 avdd.t270 27.6955
R3497 avdd.n1316 avdd.t464 27.6955
R3498 avdd.n1380 avdd.t241 27.6955
R3499 avdd.n1380 avdd.t458 27.6955
R3500 avdd.n1232 avdd.t466 27.6955
R3501 avdd.n1232 avdd.t321 27.6955
R3502 avdd.n1234 avdd.t463 27.6955
R3503 avdd.n1234 avdd.t298 27.6955
R3504 avdd.n1236 avdd.t465 27.6955
R3505 avdd.n1236 avdd.t312 27.6955
R3506 avdd.n1238 avdd.t461 27.6955
R3507 avdd.n1238 avdd.t292 27.6955
R3508 avdd.n1240 avdd.t147 27.6955
R3509 avdd.n1240 avdd.t243 27.6955
R3510 avdd.n1242 avdd.t127 27.6955
R3511 avdd.n1242 avdd.t285 27.6955
R3512 avdd.n1244 avdd.t146 27.6955
R3513 avdd.n1244 avdd.t237 27.6955
R3514 avdd.n1246 avdd.t124 27.6955
R3515 avdd.n1246 avdd.t378 27.6955
R3516 avdd.n1248 avdd.t150 27.6955
R3517 avdd.n1248 avdd.t360 27.6955
R3518 avdd.n1250 avdd.t149 27.6955
R3519 avdd.n1250 avdd.t357 27.6955
R3520 avdd.n1252 avdd.t138 27.6955
R3521 avdd.n1252 avdd.t305 27.6955
R3522 avdd.n1255 avdd.t132 27.6955
R3523 avdd.n1255 avdd.t278 27.6955
R3524 avdd.n1356 avdd.t597 27.6955
R3525 avdd.n1356 avdd.t601 27.6955
R3526 avdd.n1358 avdd.t587 27.6955
R3527 avdd.n1358 avdd.t591 27.6955
R3528 avdd.n1360 avdd.t599 27.6955
R3529 avdd.n1360 avdd.t589 27.6955
R3530 avdd.n1362 avdd.t595 27.6955
R3531 avdd.n1362 avdd.t605 27.6955
R3532 avdd.t324 avdd.n1584 26.7523
R3533 avdd.n1553 avdd.t263 25.5567
R3534 avdd.n1578 avdd.t230 25.5567
R3535 avdd.n1560 avdd.t370 25.4942
R3536 avdd.t573 avdd.t448 25.0145
R3537 avdd.n311 avdd.t161 23.5572
R3538 avdd.n283 avdd.t521 23.5572
R3539 avdd.n255 avdd.t455 23.5572
R3540 avdd.n227 avdd.t583 23.5572
R3541 avdd.n199 avdd.t407 23.5572
R3542 avdd.n171 avdd.t122 23.5572
R3543 avdd.n143 avdd.t516 23.5572
R3544 avdd.n115 avdd.t488 23.5572
R3545 avdd.n82 avdd.t53 23.5572
R3546 avdd.n647 avdd.t418 23.5572
R3547 avdd.n619 avdd.t498 23.5572
R3548 avdd.n591 avdd.t443 23.5572
R3549 avdd.n563 avdd.t537 23.5572
R3550 avdd.n535 avdd.t113 23.5572
R3551 avdd.n507 avdd.t55 23.5572
R3552 avdd.n479 avdd.t606 23.5572
R3553 avdd.n451 avdd.t11 23.5572
R3554 avdd.n418 avdd.t9 23.5572
R3555 avdd.t351 avdd.t448 22.3534
R3556 avdd.n1487 avdd.n1484 21.9177
R3557 avdd.n1499 avdd.n1498 20.3986
R3558 avdd.n1498 avdd.n1445 20.2792
R3559 avdd.n74 avdd 20.0949
R3560 avdd.n410 avdd 20.0949
R3561 avdd.n1464 avdd.n1444 19.4414
R3562 avdd.n1474 avdd.n1473 18.824
R3563 avdd.n79 avdd 18.3657
R3564 avdd.n415 avdd 18.3657
R3565 avdd.n311 avdd.t154 17.8272
R3566 avdd.n283 avdd.t518 17.8272
R3567 avdd.n255 avdd.t576 17.8272
R3568 avdd.n227 avdd.t173 17.8272
R3569 avdd.n199 avdd.t423 17.8272
R3570 avdd.n171 avdd.t1 17.8272
R3571 avdd.n143 avdd.t525 17.8272
R3572 avdd.n115 avdd.t451 17.8272
R3573 avdd.n82 avdd.t566 17.8272
R3574 avdd.n647 avdd.t216 17.8272
R3575 avdd.n619 avdd.t111 17.8272
R3576 avdd.n591 avdd.t495 17.8272
R3577 avdd.n563 avdd.t117 17.8272
R3578 avdd.n535 avdd.t538 17.8272
R3579 avdd.n507 avdd.t223 17.8272
R3580 avdd.n479 avdd.t529 17.8272
R3581 avdd.n451 avdd.t534 17.8272
R3582 avdd.n418 avdd.t222 17.8272
R3583 avdd.n1126 avdd.n1122 17.7802
R3584 avdd.n1166 avdd.n961 17.7802
R3585 avdd.n1372 avdd.n1368 17.7802
R3586 avdd.n1412 avdd.n1207 17.7802
R3587 avdd.n335 avdd.n334 17.7258
R3588 avdd.n307 avdd.n306 17.7258
R3589 avdd.n279 avdd.n278 17.7258
R3590 avdd.n251 avdd.n250 17.7258
R3591 avdd.n223 avdd.n222 17.7258
R3592 avdd.n195 avdd.n194 17.7258
R3593 avdd.n167 avdd.n166 17.7258
R3594 avdd.n139 avdd.n138 17.7258
R3595 avdd.n111 avdd.n110 17.7258
R3596 avdd.n671 avdd.n670 17.7258
R3597 avdd.n643 avdd.n642 17.7258
R3598 avdd.n615 avdd.n614 17.7258
R3599 avdd.n587 avdd.n586 17.7258
R3600 avdd.n559 avdd.n558 17.7258
R3601 avdd.n531 avdd.n530 17.7258
R3602 avdd.n503 avdd.n502 17.7258
R3603 avdd.n475 avdd.n474 17.7258
R3604 avdd.n447 avdd.n446 17.7258
R3605 avdd.n79 avdd.n78 17.3701
R3606 avdd.n78 avdd.n73 17.3701
R3607 avdd.n415 avdd.n414 17.3701
R3608 avdd.n414 avdd.n409 17.3701
R3609 avdd.n1580 avdd.n1543 16.6169
R3610 avdd.t446 avdd.t163 16.4991
R3611 avdd.n1580 avdd.n1569 16.3798
R3612 avdd.n1526 avdd.n1525 14.9605
R3613 avdd.n1533 avdd.n1532 14.9605
R3614 avdd.n1461 avdd.n1456 14.6829
R3615 avdd.n1550 avdd.n1549 14.6449
R3616 avdd.n953 avdd.t226 14.6083
R3617 avdd.n1133 avdd.t273 14.6083
R3618 avdd.n1199 avdd.t277 14.6083
R3619 avdd.n1379 avdd.t239 14.6083
R3620 avdd.n1488 avdd.n1487 14.4431
R3621 avdd.n1184 avdd.t314 14.4262
R3622 avdd.n1182 avdd.t317 14.4262
R3623 avdd.n1180 avdd.t332 14.4262
R3624 avdd.n1178 avdd.t327 14.4262
R3625 avdd.n1176 avdd.t388 14.4262
R3626 avdd.n1174 avdd.t340 14.4262
R3627 avdd.n1172 avdd.t393 14.4262
R3628 avdd.n1091 avdd.t366 14.4262
R3629 avdd.n1086 avdd.t368 14.4262
R3630 avdd.n1083 avdd.t382 14.4262
R3631 avdd.n1080 avdd.t375 14.4262
R3632 avdd.n1077 avdd.t245 14.4262
R3633 avdd.n1072 avdd.t391 14.4262
R3634 avdd.n1069 avdd.t255 14.4262
R3635 avdd.n1430 avdd.t242 14.4262
R3636 avdd.n1428 avdd.t284 14.4262
R3637 avdd.n1426 avdd.t235 14.4262
R3638 avdd.n1424 avdd.t377 14.4262
R3639 avdd.n1422 avdd.t359 14.4262
R3640 avdd.n1420 avdd.t356 14.4262
R3641 avdd.n1418 avdd.t304 14.4262
R3642 avdd.n1337 avdd.t275 14.4262
R3643 avdd.n1332 avdd.t330 14.4262
R3644 avdd.n1329 avdd.t271 14.4262
R3645 avdd.n1326 avdd.t325 14.4262
R3646 avdd.n1323 avdd.t307 14.4262
R3647 avdd.n1318 avdd.t300 14.4262
R3648 avdd.n1315 avdd.t269 14.4262
R3649 avdd.n1192 avdd.t250 14.4191
R3650 avdd.n1190 avdd.t260 14.4191
R3651 avdd.n1188 avdd.t257 14.4191
R3652 avdd.n1186 avdd.t294 14.4191
R3653 avdd.n1105 avdd.t282 14.4191
R3654 avdd.n1100 avdd.t289 14.4191
R3655 avdd.n1097 avdd.t287 14.4191
R3656 avdd.n1094 avdd.t352 14.4191
R3657 avdd.n1438 avdd.t320 14.4191
R3658 avdd.n1436 avdd.t297 14.4191
R3659 avdd.n1434 avdd.t311 14.4191
R3660 avdd.n1432 avdd.t291 14.4191
R3661 avdd.n1351 avdd.t364 14.4191
R3662 avdd.n1346 avdd.t348 14.4191
R3663 avdd.n1343 avdd.t354 14.4191
R3664 avdd.n1340 avdd.t346 14.4191
R3665 avdd.n1568 avdd.n1549 14.4078
R3666 avdd.n1586 avdd.n1585 14.2313
R3667 avdd.t324 avdd.n1586 14.2313
R3668 avdd.n1588 avdd.n1587 14.2313
R3669 avdd.n1587 avdd.t324 14.2313
R3670 avdd.n1471 avdd.n1462 14.1829
R3671 avdd.n1119 avdd.n1118 14.0622
R3672 avdd.n1365 avdd.n1364 14.0622
R3673 avdd.n1472 avdd.n674 13.9971
R3674 avdd.n1651 avdd.n1650 13.8347
R3675 avdd.n1641 avdd.n1640 13.8322
R3676 avdd.n949 avdd.n948 13.822
R3677 avdd.n1643 avdd.n950 13.822
R3678 avdd.n1171 avdd.n1170 13.8005
R3679 avdd.n1158 avdd.n1157 13.8005
R3680 avdd.n1024 avdd.n980 13.8005
R3681 avdd.n1008 avdd.n955 13.8005
R3682 avdd.n1131 avdd.n1130 13.8005
R3683 avdd.n1108 avdd.n1038 13.8005
R3684 avdd.n1417 avdd.n1416 13.8005
R3685 avdd.n1404 avdd.n1403 13.8005
R3686 avdd.n1270 avdd.n1226 13.8005
R3687 avdd.n1254 avdd.n1201 13.8005
R3688 avdd.n1377 avdd.n1376 13.8005
R3689 avdd.n1354 avdd.n1284 13.8005
R3690 avdd.n94 avdd.t565 13.7868
R3691 avdd.n430 avdd.t221 13.7868
R3692 avdd.n1023 avdd.n983 13.436
R3693 avdd.n1150 avdd.n1011 13.436
R3694 avdd.n1137 avdd.n1136 13.436
R3695 avdd.n1269 avdd.n1229 13.436
R3696 avdd.n1396 avdd.n1257 13.436
R3697 avdd.n1383 avdd.n1382 13.436
R3698 avdd.n1140 avdd.n1139 13.177
R3699 avdd.n1386 avdd.n1385 13.177
R3700 avdd.n1031 avdd.n1030 13.0943
R3701 avdd.n1030 avdd.n1029 13.0943
R3702 avdd.n1277 avdd.n1276 13.0943
R3703 avdd.n1276 avdd.n1275 13.0943
R3704 avdd.n334 avdd.n333 12.541
R3705 avdd.n306 avdd.n305 12.541
R3706 avdd.n278 avdd.n277 12.541
R3707 avdd.n250 avdd.n249 12.541
R3708 avdd.n222 avdd.n221 12.541
R3709 avdd.n194 avdd.n193 12.541
R3710 avdd.n166 avdd.n165 12.541
R3711 avdd.n138 avdd.n137 12.541
R3712 avdd.n110 avdd.n109 12.541
R3713 avdd.n670 avdd.n669 12.541
R3714 avdd.n642 avdd.n641 12.541
R3715 avdd.n614 avdd.n613 12.541
R3716 avdd.n586 avdd.n585 12.541
R3717 avdd.n558 avdd.n557 12.541
R3718 avdd.n530 avdd.n529 12.541
R3719 avdd.n502 avdd.n501 12.541
R3720 avdd.n474 avdd.n473 12.541
R3721 avdd.n446 avdd.n445 12.541
R3722 avdd.n326 avdd 12.424
R3723 avdd.n298 avdd 12.424
R3724 avdd.n270 avdd 12.424
R3725 avdd.n242 avdd 12.424
R3726 avdd.n214 avdd 12.424
R3727 avdd.n186 avdd 12.424
R3728 avdd.n158 avdd 12.424
R3729 avdd.n130 avdd 12.424
R3730 avdd.n102 avdd 12.424
R3731 avdd.n662 avdd 12.424
R3732 avdd.n634 avdd 12.424
R3733 avdd.n606 avdd 12.424
R3734 avdd.n578 avdd 12.424
R3735 avdd.n550 avdd 12.424
R3736 avdd.n522 avdd 12.424
R3737 avdd.n494 avdd 12.424
R3738 avdd.n466 avdd 12.424
R3739 avdd.n438 avdd 12.424
R3740 avdd.n1470 avdd.n1460 11.2946
R3741 avdd.n1484 avdd.n1445 11.1593
R3742 avdd.n1548 avdd.n1547 11.0005
R3743 avdd.n1582 avdd.n1581 11.0005
R3744 avdd.n1031 avdd.n977 10.9402
R3745 avdd.n1029 avdd.n977 10.9402
R3746 avdd.n1277 avdd.n1223 10.9402
R3747 avdd.n1275 avdd.n1223 10.9402
R3748 avdd.n1634 avdd.n1633 10.8829
R3749 avdd.n1631 avdd.n1626 10.8829
R3750 avdd.n1646 avdd.n1645 10.8829
R3751 avdd.n1648 avdd.n1647 10.8829
R3752 avdd.n1535 avdd.n1534 10.2783
R3753 avdd.n1537 avdd.n1536 10.2783
R3754 avdd.n1538 avdd.n1537 10.2783
R3755 avdd.n1516 avdd.n1513 10.2783
R3756 avdd.n1517 avdd.n1516 10.2783
R3757 avdd.n1511 avdd.n1508 10.2783
R3758 avdd.n1544 avdd.n1511 10.2783
R3759 avdd.n1547 avdd.n1546 10.2783
R3760 avdd.n1583 avdd.n1582 10.2783
R3761 avdd.n1584 avdd.n1583 10.2783
R3762 avdd.t421 avdd.t50 10.0269
R3763 avdd.t102 avdd.t6 10.0269
R3764 avdd.n1153 avdd.n984 9.71534
R3765 avdd.n1399 avdd.n1230 9.71534
R3766 avdd.n331 avdd.n330 9.5406
R3767 avdd.n303 avdd.n302 9.5406
R3768 avdd.n275 avdd.n274 9.5406
R3769 avdd.n247 avdd.n246 9.5406
R3770 avdd.n219 avdd.n218 9.5406
R3771 avdd.n191 avdd.n190 9.5406
R3772 avdd.n163 avdd.n162 9.5406
R3773 avdd.n135 avdd.n134 9.5406
R3774 avdd.n107 avdd.n106 9.5406
R3775 avdd.n667 avdd.n666 9.5406
R3776 avdd.n639 avdd.n638 9.5406
R3777 avdd.n611 avdd.n610 9.5406
R3778 avdd.n583 avdd.n582 9.5406
R3779 avdd.n555 avdd.n554 9.5406
R3780 avdd.n527 avdd.n526 9.5406
R3781 avdd.n499 avdd.n498 9.5406
R3782 avdd.n471 avdd.n470 9.5406
R3783 avdd.n443 avdd.n442 9.5406
R3784 avdd.n1455 avdd.n674 9.42955
R3785 avdd.n1481 avdd.n1480 9.41227
R3786 avdd.n80 avdd.n73 9.3005
R3787 avdd.n108 avdd.n107 9.3005
R3788 avdd.n107 avdd.n105 9.3005
R3789 avdd.n136 avdd.n135 9.3005
R3790 avdd.n135 avdd.n133 9.3005
R3791 avdd.n164 avdd.n163 9.3005
R3792 avdd.n163 avdd.n161 9.3005
R3793 avdd.n192 avdd.n191 9.3005
R3794 avdd.n191 avdd.n189 9.3005
R3795 avdd.n220 avdd.n219 9.3005
R3796 avdd.n219 avdd.n217 9.3005
R3797 avdd.n248 avdd.n247 9.3005
R3798 avdd.n247 avdd.n245 9.3005
R3799 avdd.n276 avdd.n275 9.3005
R3800 avdd.n275 avdd.n273 9.3005
R3801 avdd.n304 avdd.n303 9.3005
R3802 avdd.n303 avdd.n301 9.3005
R3803 avdd.n332 avdd.n331 9.3005
R3804 avdd.n331 avdd.n329 9.3005
R3805 avdd.n80 avdd.n79 9.3005
R3806 avdd.n87 avdd.n86 9.3005
R3807 avdd.n88 avdd.n87 9.3005
R3808 avdd.n119 avdd.n118 9.3005
R3809 avdd.n118 avdd.n117 9.3005
R3810 avdd.n147 avdd.n146 9.3005
R3811 avdd.n146 avdd.n145 9.3005
R3812 avdd.n175 avdd.n174 9.3005
R3813 avdd.n174 avdd.n173 9.3005
R3814 avdd.n203 avdd.n202 9.3005
R3815 avdd.n202 avdd.n201 9.3005
R3816 avdd.n231 avdd.n230 9.3005
R3817 avdd.n230 avdd.n229 9.3005
R3818 avdd.n259 avdd.n258 9.3005
R3819 avdd.n258 avdd.n257 9.3005
R3820 avdd.n287 avdd.n286 9.3005
R3821 avdd.n286 avdd.n285 9.3005
R3822 avdd.n315 avdd.n314 9.3005
R3823 avdd.n314 avdd.n313 9.3005
R3824 avdd.n77 avdd.n76 9.3005
R3825 avdd.n81 avdd.n71 9.3005
R3826 avdd.n91 avdd.n90 9.3005
R3827 avdd.n89 avdd.n72 9.3005
R3828 avdd.n84 avdd.n68 9.3005
R3829 avdd.n85 avdd.n65 9.3005
R3830 avdd.n104 avdd.n103 9.3005
R3831 avdd.n102 avdd.n64 9.3005
R3832 avdd.n126 avdd.n125 9.3005
R3833 avdd.n124 avdd.n63 9.3005
R3834 avdd.n123 avdd.n122 9.3005
R3835 avdd.n121 avdd.n120 9.3005
R3836 avdd.n114 avdd.n57 9.3005
R3837 avdd.n132 avdd.n131 9.3005
R3838 avdd.n130 avdd.n56 9.3005
R3839 avdd.n154 avdd.n153 9.3005
R3840 avdd.n152 avdd.n55 9.3005
R3841 avdd.n151 avdd.n150 9.3005
R3842 avdd.n149 avdd.n148 9.3005
R3843 avdd.n142 avdd.n49 9.3005
R3844 avdd.n160 avdd.n159 9.3005
R3845 avdd.n158 avdd.n48 9.3005
R3846 avdd.n182 avdd.n181 9.3005
R3847 avdd.n180 avdd.n47 9.3005
R3848 avdd.n179 avdd.n178 9.3005
R3849 avdd.n177 avdd.n176 9.3005
R3850 avdd.n170 avdd.n41 9.3005
R3851 avdd.n188 avdd.n187 9.3005
R3852 avdd.n186 avdd.n40 9.3005
R3853 avdd.n210 avdd.n209 9.3005
R3854 avdd.n208 avdd.n39 9.3005
R3855 avdd.n207 avdd.n206 9.3005
R3856 avdd.n205 avdd.n204 9.3005
R3857 avdd.n198 avdd.n33 9.3005
R3858 avdd.n216 avdd.n215 9.3005
R3859 avdd.n214 avdd.n32 9.3005
R3860 avdd.n238 avdd.n237 9.3005
R3861 avdd.n236 avdd.n31 9.3005
R3862 avdd.n235 avdd.n234 9.3005
R3863 avdd.n233 avdd.n232 9.3005
R3864 avdd.n226 avdd.n25 9.3005
R3865 avdd.n244 avdd.n243 9.3005
R3866 avdd.n242 avdd.n24 9.3005
R3867 avdd.n266 avdd.n265 9.3005
R3868 avdd.n264 avdd.n23 9.3005
R3869 avdd.n263 avdd.n262 9.3005
R3870 avdd.n261 avdd.n260 9.3005
R3871 avdd.n254 avdd.n17 9.3005
R3872 avdd.n272 avdd.n271 9.3005
R3873 avdd.n270 avdd.n16 9.3005
R3874 avdd.n294 avdd.n293 9.3005
R3875 avdd.n292 avdd.n15 9.3005
R3876 avdd.n291 avdd.n290 9.3005
R3877 avdd.n289 avdd.n288 9.3005
R3878 avdd.n282 avdd.n9 9.3005
R3879 avdd.n300 avdd.n299 9.3005
R3880 avdd.n298 avdd.n8 9.3005
R3881 avdd.n322 avdd.n321 9.3005
R3882 avdd.n320 avdd.n7 9.3005
R3883 avdd.n319 avdd.n318 9.3005
R3884 avdd.n317 avdd.n316 9.3005
R3885 avdd.n310 avdd.n1 9.3005
R3886 avdd.n328 avdd.n327 9.3005
R3887 avdd.n326 avdd.n0 9.3005
R3888 avdd.n416 avdd.n409 9.3005
R3889 avdd.n444 avdd.n443 9.3005
R3890 avdd.n443 avdd.n441 9.3005
R3891 avdd.n472 avdd.n471 9.3005
R3892 avdd.n471 avdd.n469 9.3005
R3893 avdd.n500 avdd.n499 9.3005
R3894 avdd.n499 avdd.n497 9.3005
R3895 avdd.n528 avdd.n527 9.3005
R3896 avdd.n527 avdd.n525 9.3005
R3897 avdd.n556 avdd.n555 9.3005
R3898 avdd.n555 avdd.n553 9.3005
R3899 avdd.n584 avdd.n583 9.3005
R3900 avdd.n583 avdd.n581 9.3005
R3901 avdd.n612 avdd.n611 9.3005
R3902 avdd.n611 avdd.n609 9.3005
R3903 avdd.n640 avdd.n639 9.3005
R3904 avdd.n639 avdd.n637 9.3005
R3905 avdd.n668 avdd.n667 9.3005
R3906 avdd.n667 avdd.n665 9.3005
R3907 avdd.n416 avdd.n415 9.3005
R3908 avdd.n423 avdd.n422 9.3005
R3909 avdd.n424 avdd.n423 9.3005
R3910 avdd.n455 avdd.n454 9.3005
R3911 avdd.n454 avdd.n453 9.3005
R3912 avdd.n483 avdd.n482 9.3005
R3913 avdd.n482 avdd.n481 9.3005
R3914 avdd.n511 avdd.n510 9.3005
R3915 avdd.n510 avdd.n509 9.3005
R3916 avdd.n539 avdd.n538 9.3005
R3917 avdd.n538 avdd.n537 9.3005
R3918 avdd.n567 avdd.n566 9.3005
R3919 avdd.n566 avdd.n565 9.3005
R3920 avdd.n595 avdd.n594 9.3005
R3921 avdd.n594 avdd.n593 9.3005
R3922 avdd.n623 avdd.n622 9.3005
R3923 avdd.n622 avdd.n621 9.3005
R3924 avdd.n651 avdd.n650 9.3005
R3925 avdd.n650 avdd.n649 9.3005
R3926 avdd.n413 avdd.n412 9.3005
R3927 avdd.n417 avdd.n407 9.3005
R3928 avdd.n427 avdd.n426 9.3005
R3929 avdd.n425 avdd.n408 9.3005
R3930 avdd.n420 avdd.n404 9.3005
R3931 avdd.n421 avdd.n401 9.3005
R3932 avdd.n440 avdd.n439 9.3005
R3933 avdd.n438 avdd.n400 9.3005
R3934 avdd.n462 avdd.n461 9.3005
R3935 avdd.n460 avdd.n399 9.3005
R3936 avdd.n459 avdd.n458 9.3005
R3937 avdd.n457 avdd.n456 9.3005
R3938 avdd.n450 avdd.n393 9.3005
R3939 avdd.n468 avdd.n467 9.3005
R3940 avdd.n466 avdd.n392 9.3005
R3941 avdd.n490 avdd.n489 9.3005
R3942 avdd.n488 avdd.n391 9.3005
R3943 avdd.n487 avdd.n486 9.3005
R3944 avdd.n485 avdd.n484 9.3005
R3945 avdd.n478 avdd.n385 9.3005
R3946 avdd.n496 avdd.n495 9.3005
R3947 avdd.n494 avdd.n384 9.3005
R3948 avdd.n518 avdd.n517 9.3005
R3949 avdd.n516 avdd.n383 9.3005
R3950 avdd.n515 avdd.n514 9.3005
R3951 avdd.n513 avdd.n512 9.3005
R3952 avdd.n506 avdd.n377 9.3005
R3953 avdd.n524 avdd.n523 9.3005
R3954 avdd.n522 avdd.n376 9.3005
R3955 avdd.n546 avdd.n545 9.3005
R3956 avdd.n544 avdd.n375 9.3005
R3957 avdd.n543 avdd.n542 9.3005
R3958 avdd.n541 avdd.n540 9.3005
R3959 avdd.n534 avdd.n369 9.3005
R3960 avdd.n552 avdd.n551 9.3005
R3961 avdd.n550 avdd.n368 9.3005
R3962 avdd.n574 avdd.n573 9.3005
R3963 avdd.n572 avdd.n367 9.3005
R3964 avdd.n571 avdd.n570 9.3005
R3965 avdd.n569 avdd.n568 9.3005
R3966 avdd.n562 avdd.n361 9.3005
R3967 avdd.n580 avdd.n579 9.3005
R3968 avdd.n578 avdd.n360 9.3005
R3969 avdd.n602 avdd.n601 9.3005
R3970 avdd.n600 avdd.n359 9.3005
R3971 avdd.n599 avdd.n598 9.3005
R3972 avdd.n597 avdd.n596 9.3005
R3973 avdd.n590 avdd.n353 9.3005
R3974 avdd.n608 avdd.n607 9.3005
R3975 avdd.n606 avdd.n352 9.3005
R3976 avdd.n630 avdd.n629 9.3005
R3977 avdd.n628 avdd.n351 9.3005
R3978 avdd.n627 avdd.n626 9.3005
R3979 avdd.n625 avdd.n624 9.3005
R3980 avdd.n618 avdd.n345 9.3005
R3981 avdd.n636 avdd.n635 9.3005
R3982 avdd.n634 avdd.n344 9.3005
R3983 avdd.n658 avdd.n657 9.3005
R3984 avdd.n656 avdd.n343 9.3005
R3985 avdd.n655 avdd.n654 9.3005
R3986 avdd.n653 avdd.n652 9.3005
R3987 avdd.n646 avdd.n337 9.3005
R3988 avdd.n664 avdd.n663 9.3005
R3989 avdd.n662 avdd.n336 9.3005
R3990 avdd.n1628 avdd.n1625 9.3005
R3991 avdd.n1637 avdd.n1609 9.3005
R3992 avdd.n686 avdd.n685 9.3005
R3993 avdd.n687 avdd.n686 9.3005
R3994 avdd.n677 avdd.n675 9.3005
R3995 avdd.n684 avdd.n683 9.3005
R3996 avdd.n682 avdd.n676 9.3005
R3997 avdd.n1602 avdd.n1601 9.3005
R3998 avdd.n1581 avdd.n1580 9.3005
R3999 avdd.n1549 avdd.n1548 9.3005
R4000 avdd.n1644 avdd.n1643 9.3005
R4001 avdd.n1641 avdd.n691 9.3005
R4002 avdd.n1650 avdd.n1649 9.3005
R4003 avdd.n948 avdd.n694 9.3005
R4004 avdd.n926 avdd.n700 9.3005
R4005 avdd.n927 avdd.n926 9.3005
R4006 avdd.n915 avdd.n707 9.3005
R4007 avdd.n916 avdd.n915 9.3005
R4008 avdd.n715 avdd.n714 9.3005
R4009 avdd.n716 avdd.n715 9.3005
R4010 avdd.n903 avdd.n902 9.3005
R4011 avdd.n902 avdd.n901 9.3005
R4012 avdd.n890 avdd.n727 9.3005
R4013 avdd.n891 avdd.n890 9.3005
R4014 avdd.n735 avdd.n734 9.3005
R4015 avdd.n736 avdd.n735 9.3005
R4016 avdd.n878 avdd.n877 9.3005
R4017 avdd.n877 avdd.n876 9.3005
R4018 avdd.n865 avdd.n747 9.3005
R4019 avdd.n866 avdd.n865 9.3005
R4020 avdd.n755 avdd.n754 9.3005
R4021 avdd.n756 avdd.n755 9.3005
R4022 avdd.n853 avdd.n852 9.3005
R4023 avdd.n852 avdd.n851 9.3005
R4024 avdd.n840 avdd.n767 9.3005
R4025 avdd.n841 avdd.n840 9.3005
R4026 avdd.n775 avdd.n774 9.3005
R4027 avdd.n776 avdd.n775 9.3005
R4028 avdd.n828 avdd.n827 9.3005
R4029 avdd.n827 avdd.n826 9.3005
R4030 avdd.n815 avdd.n787 9.3005
R4031 avdd.n816 avdd.n815 9.3005
R4032 avdd.n795 avdd.n794 9.3005
R4033 avdd.n796 avdd.n795 9.3005
R4034 avdd.n803 avdd.n802 9.3005
R4035 avdd.n802 avdd.n801 9.3005
R4036 avdd.n932 avdd.n931 9.3005
R4037 avdd.n930 avdd.n696 9.3005
R4038 avdd.n929 avdd.n928 9.3005
R4039 avdd.n925 avdd.n924 9.3005
R4040 avdd.n702 avdd.n701 9.3005
R4041 avdd.n918 avdd.n917 9.3005
R4042 avdd.n914 avdd.n913 9.3005
R4043 avdd.n709 avdd.n708 9.3005
R4044 avdd.n713 avdd.n712 9.3005
R4045 avdd.n906 avdd.n717 9.3005
R4046 avdd.n905 avdd.n904 9.3005
R4047 avdd.n719 avdd.n718 9.3005
R4048 avdd.n900 avdd.n899 9.3005
R4049 avdd.n721 avdd.n720 9.3005
R4050 avdd.n893 avdd.n892 9.3005
R4051 avdd.n889 avdd.n888 9.3005
R4052 avdd.n729 avdd.n728 9.3005
R4053 avdd.n733 avdd.n732 9.3005
R4054 avdd.n881 avdd.n737 9.3005
R4055 avdd.n880 avdd.n879 9.3005
R4056 avdd.n739 avdd.n738 9.3005
R4057 avdd.n875 avdd.n874 9.3005
R4058 avdd.n741 avdd.n740 9.3005
R4059 avdd.n868 avdd.n867 9.3005
R4060 avdd.n864 avdd.n863 9.3005
R4061 avdd.n749 avdd.n748 9.3005
R4062 avdd.n753 avdd.n752 9.3005
R4063 avdd.n856 avdd.n757 9.3005
R4064 avdd.n855 avdd.n854 9.3005
R4065 avdd.n759 avdd.n758 9.3005
R4066 avdd.n850 avdd.n849 9.3005
R4067 avdd.n761 avdd.n760 9.3005
R4068 avdd.n843 avdd.n842 9.3005
R4069 avdd.n839 avdd.n838 9.3005
R4070 avdd.n769 avdd.n768 9.3005
R4071 avdd.n773 avdd.n772 9.3005
R4072 avdd.n831 avdd.n777 9.3005
R4073 avdd.n830 avdd.n829 9.3005
R4074 avdd.n779 avdd.n778 9.3005
R4075 avdd.n825 avdd.n824 9.3005
R4076 avdd.n781 avdd.n780 9.3005
R4077 avdd.n818 avdd.n817 9.3005
R4078 avdd.n814 avdd.n813 9.3005
R4079 avdd.n789 avdd.n788 9.3005
R4080 avdd.n793 avdd.n792 9.3005
R4081 avdd.n806 avdd.n797 9.3005
R4082 avdd.n805 avdd.n804 9.3005
R4083 avdd.n800 avdd.n799 9.3005
R4084 avdd.n1501 avdd.n1500 9.27144
R4085 avdd.n1642 avdd.n1641 9.2699
R4086 avdd.n1643 avdd.n1642 9.2699
R4087 avdd.n1472 avdd.n1471 8.94982
R4088 avdd.n967 avdd.n965 8.40959
R4089 avdd.n967 avdd.n961 8.40959
R4090 avdd.n971 avdd.n966 8.40959
R4091 avdd.n971 avdd.n961 8.40959
R4092 avdd.n1125 avdd.n1124 8.40959
R4093 avdd.n1126 avdd.n1125 8.40959
R4094 avdd.n1165 avdd.n1164 8.40959
R4095 avdd.n1166 avdd.n1165 8.40959
R4096 avdd.n1213 avdd.n1211 8.40959
R4097 avdd.n1213 avdd.n1207 8.40959
R4098 avdd.n1217 avdd.n1212 8.40959
R4099 avdd.n1217 avdd.n1207 8.40959
R4100 avdd.n1371 avdd.n1370 8.40959
R4101 avdd.n1372 avdd.n1371 8.40959
R4102 avdd.n1411 avdd.n1410 8.40959
R4103 avdd.n1412 avdd.n1411 8.40959
R4104 avdd.n1138 avdd.n1021 8.24855
R4105 avdd.n1384 avdd.n1267 8.24855
R4106 avdd.n1197 avdd.n1196 8.24253
R4107 avdd.n1443 avdd.n1442 8.24253
R4108 avdd.n1148 avdd.n1011 8.18605
R4109 avdd.n1394 avdd.n1257 8.18605
R4110 avdd.n1149 avdd.n1148 8.17238
R4111 avdd.n1395 avdd.n1394 8.17238
R4112 avdd.n1138 avdd.n1137 8.10988
R4113 avdd.n1384 avdd.n1383 8.10988
R4114 avdd.n1606 avdd.n1605 7.90948
R4115 avdd.n1108 avdd.n1107 7.90079
R4116 avdd.n1354 avdd.n1353 7.90079
R4117 avdd.n1602 avdd.n1506 7.55653
R4118 avdd.n1519 avdd.n1506 7.55653
R4119 avdd.n1598 avdd.n1597 7.4005
R4120 avdd.t351 avdd.n1598 7.4005
R4121 avdd.n1600 avdd.n1599 7.4005
R4122 avdd.n1599 avdd.t351 7.4005
R4123 avdd.n1022 avdd.n1011 7.29542
R4124 avdd.n1268 avdd.n1257 7.29542
R4125 avdd.n1606 avdd.n950 7.06613
R4126 avdd.n1519 avdd.n1507 7.06516
R4127 avdd.n1602 avdd.n1507 7.06516
R4128 avdd.n330 avdd 7.01471
R4129 avdd.n302 avdd 7.01471
R4130 avdd.n274 avdd 7.01471
R4131 avdd.n246 avdd 7.01471
R4132 avdd.n218 avdd 7.01471
R4133 avdd.n190 avdd 7.01471
R4134 avdd.n162 avdd 7.01471
R4135 avdd.n134 avdd 7.01471
R4136 avdd.n106 avdd 7.01471
R4137 avdd.n666 avdd 7.01471
R4138 avdd.n638 avdd 7.01471
R4139 avdd.n610 avdd 7.01471
R4140 avdd.n582 avdd 7.01471
R4141 avdd.n554 avdd 7.01471
R4142 avdd.n526 avdd 7.01471
R4143 avdd.n498 avdd 7.01471
R4144 avdd.n470 avdd 7.01471
R4145 avdd.n442 avdd 7.01471
R4146 avdd.n1137 avdd.n1023 6.77003
R4147 avdd.n1021 avdd.n1020 6.77003
R4148 avdd.n1383 avdd.n1269 6.77003
R4149 avdd.n1267 avdd.n1266 6.77003
R4150 avdd.n1040 avdd.n1035 6.60764
R4151 avdd.n1122 avdd.n1035 6.60764
R4152 avdd.n1121 avdd.n1120 6.60764
R4153 avdd.n1122 avdd.n1121 6.60764
R4154 avdd.n1286 avdd.n1281 6.60764
R4155 avdd.n1368 avdd.n1281 6.60764
R4156 avdd.n1367 avdd.n1366 6.60764
R4157 avdd.n1368 avdd.n1367 6.60764
R4158 avdd.n1149 avdd.n1012 6.59816
R4159 avdd.n1395 avdd.n1258 6.59816
R4160 avdd.n1153 avdd.n1152 6.47706
R4161 avdd.n1399 avdd.n1398 6.47706
R4162 avdd.n1639 avdd.n1638 5.7183
R4163 avdd.n1554 avdd.n1553 5.70732
R4164 avdd.n1579 avdd.n1578 5.70732
R4165 avdd.n1561 avdd.n1560 5.70732
R4166 avdd.n1554 avdd.n1549 5.70369
R4167 avdd.n1625 avdd.n1624 5.70305
R4168 avdd.n1580 avdd.n1579 5.70274
R4169 avdd.n1520 avdd.n1519 5.70242
R4170 avdd.n1638 avdd.n1637 5.6605
R4171 avdd.n1603 avdd.n1602 5.6605
R4172 avdd.n1566 avdd.n1565 5.6605
R4173 avdd.n1622 avdd.t83 5.5395
R4174 avdd.n1622 avdd.t65 5.5395
R4175 avdd.n1620 avdd.t87 5.5395
R4176 avdd.n1620 avdd.t67 5.5395
R4177 avdd.n1618 avdd.t75 5.5395
R4178 avdd.n1618 avdd.t71 5.5395
R4179 avdd.n1616 avdd.t77 5.5395
R4180 avdd.n1616 avdd.t61 5.5395
R4181 avdd.n1614 avdd.t81 5.5395
R4182 avdd.n1614 avdd.t63 5.5395
R4183 avdd.n1612 avdd.t69 5.5395
R4184 avdd.n1612 avdd.t85 5.5395
R4185 avdd.n1610 avdd.t73 5.5395
R4186 avdd.n1610 avdd.t89 5.5395
R4187 avdd.n1562 avdd.t99 5.5395
R4188 avdd.t337 avdd.n1562 5.5395
R4189 avdd.n1504 avdd.t345 5.5395
R4190 avdd.n1504 avdd.t572 5.5395
R4191 avdd.n1528 avdd.t546 5.5395
R4192 avdd.n1528 avdd.t556 5.5395
R4193 avdd.n1530 avdd.t558 5.5395
R4194 avdd.n1530 avdd.t219 5.5395
R4195 avdd.n1559 avdd.t508 5.5395
R4196 avdd.n1559 avdd.t372 5.5395
R4197 avdd.n1555 avdd.t512 5.5395
R4198 avdd.n1555 avdd.t265 5.5395
R4199 avdd.t372 avdd.n1558 5.5395
R4200 avdd.n1558 avdd.t510 5.5395
R4201 avdd.n1563 avdd.t337 5.5395
R4202 avdd.n1563 avdd.t506 5.5395
R4203 avdd.n1570 avdd.t91 5.5395
R4204 avdd.n1570 avdd.t93 5.5395
R4205 avdd.n1572 avdd.t449 5.5395
R4206 avdd.n1572 avdd.t95 5.5395
R4207 avdd.n1574 avdd.t97 5.5395
R4208 avdd.n1574 avdd.t447 5.5395
R4209 avdd.t232 avdd.n1577 5.5395
R4210 avdd.n1577 avdd.t101 5.5395
R4211 avdd.n1636 avdd.n1625 5.48326
R4212 avdd.n1637 avdd.n1636 5.48326
R4213 avdd.n704 avdd.t563 5.48127
R4214 avdd.t530 avdd.n921 5.48127
R4215 avdd.n910 avdd.t46 5.48127
R4216 avdd.n723 avdd.t408 5.48127
R4217 avdd.t104 avdd.n896 5.48127
R4218 avdd.n885 avdd.t157 5.48127
R4219 avdd.n743 avdd.t577 5.48127
R4220 avdd.t539 avdd.n871 5.48127
R4221 avdd.n860 avdd.t609 5.48127
R4222 avdd.n763 avdd.t207 5.48127
R4223 avdd.t118 avdd.n846 5.48127
R4224 avdd.n835 avdd.t579 5.48127
R4225 avdd.n783 avdd.t581 5.48127
R4226 avdd.t106 avdd.n821 5.48127
R4227 avdd.n810 avdd.t211 5.48127
R4228 avdd.n1594 avdd.n1593 5.28621
R4229 avdd.n1593 avdd.t545 5.28621
R4230 avdd.n1592 avdd.n1591 5.28621
R4231 avdd.t545 avdd.n1592 5.28621
R4232 avdd.n985 avdd.n954 5.22511
R4233 avdd.n1132 avdd.n984 5.22511
R4234 avdd.n1231 avdd.n1200 5.22511
R4235 avdd.n1378 avdd.n1230 5.22511
R4236 avdd.n1136 avdd.n1135 5.11573
R4237 avdd.n1382 avdd.n1381 5.11573
R4238 avdd.n1032 avdd.n984 4.98102
R4239 avdd.n1278 avdd.n1230 4.98102
R4240 avdd.n1028 avdd.n985 4.94972
R4241 avdd.n1274 avdd.n1231 4.94972
R4242 avdd.n1469 avdd.n1466 4.89462
R4243 avdd.n1465 avdd.n1463 4.89462
R4244 avdd.n1123 avdd.n1034 4.86892
R4245 avdd.n1126 avdd.n1123 4.86892
R4246 avdd.n1026 avdd.n960 4.86892
R4247 avdd.n1166 avdd.n960 4.86892
R4248 avdd.n1369 avdd.n1280 4.86892
R4249 avdd.n1372 avdd.n1369 4.86892
R4250 avdd.n1272 avdd.n1206 4.86892
R4251 avdd.n1412 avdd.n1206 4.86892
R4252 avdd.n673 avdd.n672 4.7853
R4253 avdd.n954 avdd.n953 4.66083
R4254 avdd.n1133 avdd.n1132 4.66083
R4255 avdd.n1200 avdd.n1199 4.66083
R4256 avdd.n1379 avdd.n1378 4.66083
R4257 avdd.n1173 avdd.n1172 4.5005
R4258 avdd.n1175 avdd.n1174 4.5005
R4259 avdd.n1177 avdd.n1176 4.5005
R4260 avdd.n1179 avdd.n1178 4.5005
R4261 avdd.n1181 avdd.n1180 4.5005
R4262 avdd.n1183 avdd.n1182 4.5005
R4263 avdd.n1185 avdd.n1184 4.5005
R4264 avdd.n1187 avdd.n1186 4.5005
R4265 avdd.n1189 avdd.n1188 4.5005
R4266 avdd.n1191 avdd.n1190 4.5005
R4267 avdd.n1193 avdd.n1192 4.5005
R4268 avdd.n1150 avdd.n1149 4.5005
R4269 avdd.n1020 avdd.n983 4.5005
R4270 avdd.n1136 avdd.n1021 4.5005
R4271 avdd.n1069 avdd.n1025 4.5005
R4272 avdd.n1072 avdd.n1068 4.5005
R4273 avdd.n1078 avdd.n1077 4.5005
R4274 avdd.n1081 avdd.n1080 4.5005
R4275 avdd.n1083 avdd.n1082 4.5005
R4276 avdd.n1086 avdd.n1066 4.5005
R4277 avdd.n1092 avdd.n1091 4.5005
R4278 avdd.n1095 avdd.n1094 4.5005
R4279 avdd.n1097 avdd.n1096 4.5005
R4280 avdd.n1100 avdd.n1064 4.5005
R4281 avdd.n1106 avdd.n1105 4.5005
R4282 avdd.n1154 avdd.n1153 4.5005
R4283 avdd.n1152 avdd.n1151 4.5005
R4284 avdd.n1419 avdd.n1418 4.5005
R4285 avdd.n1421 avdd.n1420 4.5005
R4286 avdd.n1423 avdd.n1422 4.5005
R4287 avdd.n1425 avdd.n1424 4.5005
R4288 avdd.n1427 avdd.n1426 4.5005
R4289 avdd.n1429 avdd.n1428 4.5005
R4290 avdd.n1431 avdd.n1430 4.5005
R4291 avdd.n1433 avdd.n1432 4.5005
R4292 avdd.n1435 avdd.n1434 4.5005
R4293 avdd.n1437 avdd.n1436 4.5005
R4294 avdd.n1439 avdd.n1438 4.5005
R4295 avdd.n1396 avdd.n1395 4.5005
R4296 avdd.n1266 avdd.n1229 4.5005
R4297 avdd.n1382 avdd.n1267 4.5005
R4298 avdd.n1315 avdd.n1271 4.5005
R4299 avdd.n1318 avdd.n1314 4.5005
R4300 avdd.n1324 avdd.n1323 4.5005
R4301 avdd.n1327 avdd.n1326 4.5005
R4302 avdd.n1329 avdd.n1328 4.5005
R4303 avdd.n1332 avdd.n1312 4.5005
R4304 avdd.n1338 avdd.n1337 4.5005
R4305 avdd.n1341 avdd.n1340 4.5005
R4306 avdd.n1343 avdd.n1342 4.5005
R4307 avdd.n1346 avdd.n1310 4.5005
R4308 avdd.n1352 avdd.n1351 4.5005
R4309 avdd.n1400 avdd.n1399 4.5005
R4310 avdd.n1398 avdd.n1397 4.5005
R4311 avdd.n1605 avdd.n1502 4.4965
R4312 avdd.n79 avdd 4.46111
R4313 avdd.n79 avdd 4.46111
R4314 avdd.n415 avdd 4.46111
R4315 avdd.n415 avdd 4.46111
R4316 avdd.n1194 avdd.n1193 4.45347
R4317 avdd.n1062 avdd.n1061 4.45347
R4318 avdd.n1103 avdd.n1063 4.45347
R4319 avdd.n987 avdd.n952 4.45347
R4320 avdd.n1107 avdd.n1106 4.45347
R4321 avdd.n1440 avdd.n1439 4.45347
R4322 avdd.n1308 avdd.n1307 4.45347
R4323 avdd.n1349 avdd.n1309 4.45347
R4324 avdd.n1233 avdd.n1198 4.45347
R4325 avdd.n1353 avdd.n1352 4.45347
R4326 avdd.n1151 avdd.n1150 4.39112
R4327 avdd.n1397 avdd.n1396 4.39112
R4328 avdd.n1635 avdd.n1627 4.20505
R4329 avdd.n1632 avdd.n1627 4.20505
R4330 avdd.n1630 avdd.n1629 4.20505
R4331 avdd.n1632 avdd.n1630 4.20505
R4332 avdd.n1154 avdd.n983 4.16066
R4333 avdd.n1400 avdd.n1229 4.16066
R4334 avdd.n1605 avdd.n1604 4.15861
R4335 avdd.n1490 avdd.n1489 4.14168
R4336 avdd.n1604 avdd.n1603 4.01324
R4337 avdd.n1637 avdd.n1608 3.91429
R4338 avdd.n1625 avdd.n1608 3.91429
R4339 avdd.n312 avdd 3.7406
R4340 avdd.n284 avdd 3.7406
R4341 avdd.n256 avdd 3.7406
R4342 avdd.n228 avdd 3.7406
R4343 avdd.n200 avdd 3.7406
R4344 avdd.n172 avdd 3.7406
R4345 avdd.n144 avdd 3.7406
R4346 avdd.n116 avdd 3.7406
R4347 avdd.n83 avdd 3.7406
R4348 avdd.n648 avdd 3.7406
R4349 avdd.n620 avdd 3.7406
R4350 avdd.n592 avdd 3.7406
R4351 avdd.n564 avdd 3.7406
R4352 avdd.n536 avdd 3.7406
R4353 avdd.n508 avdd 3.7406
R4354 avdd.n480 avdd 3.7406
R4355 avdd.n452 avdd 3.7406
R4356 avdd.n419 avdd 3.7406
R4357 avdd.n1460 avdd.n1459 3.55819
R4358 avdd.n1459 avdd.n1458 3.55819
R4359 avdd.n1152 avdd.n985 3.23878
R4360 avdd.n1398 avdd.n1231 3.23878
R4361 avdd.n1491 avdd.n1490 2.93701
R4362 avdd.n1492 avdd.n1491 2.93701
R4363 avdd.n1141 avdd.n1140 2.80353
R4364 avdd.n1142 avdd.n1141 2.80353
R4365 avdd.n1146 avdd.n1145 2.80353
R4366 avdd.n1145 avdd.n1144 2.80353
R4367 avdd.n1387 avdd.n1386 2.80353
R4368 avdd.n1388 avdd.n1387 2.80353
R4369 avdd.n1392 avdd.n1391 2.80353
R4370 avdd.n1391 avdd.n1390 2.80353
R4371 avdd.n672 avdd 2.67636
R4372 avdd.n1475 avdd.n1474 2.28445
R4373 avdd.n1476 avdd.n1475 2.28445
R4374 avdd.n1500 avdd.n1499 2.27397
R4375 avdd.n1604 avdd.n1503 1.97988
R4376 avdd.n1550 avdd.n1543 1.97248
R4377 avdd.n1569 avdd.n1568 1.97248
R4378 avdd.t94 avdd.n1544 1.86325
R4379 avdd.n1501 avdd 1.67975
R4380 avdd.n1029 avdd.n1028 1.61378
R4381 avdd.n1275 avdd.n1274 1.61378
R4382 avdd.n1032 avdd.n1031 1.55875
R4383 avdd.n1278 avdd.n1277 1.55875
R4384 avdd.n1446 avdd.n1444 1.5505
R4385 avdd.n1552 avdd.n1551 1.52433
R4386 avdd.n1147 avdd.n1146 1.50638
R4387 avdd.n1393 avdd.n1392 1.50638
R4388 avdd.n692 avdd.n690 1.4805
R4389 avdd.t387 avdd.n692 1.4805
R4390 avdd.n695 avdd.n693 1.4805
R4391 avdd.t387 avdd.n693 1.4805
R4392 avdd.n1567 avdd.n1566 1.31832
R4393 avdd.n948 avdd.n947 1.28283
R4394 avdd.n964 avdd.n962 1.2505
R4395 avdd.n1160 avdd.n962 1.2505
R4396 avdd.n1162 avdd.n1161 1.2505
R4397 avdd.n1161 avdd.n1160 1.2505
R4398 avdd.n1159 avdd.n1158 1.2505
R4399 avdd.n1160 avdd.n1159 1.2505
R4400 avdd.n959 avdd.n957 1.2505
R4401 avdd.n1160 avdd.n959 1.2505
R4402 avdd.n1210 avdd.n1208 1.2505
R4403 avdd.n1406 avdd.n1208 1.2505
R4404 avdd.n1408 avdd.n1407 1.2505
R4405 avdd.n1407 avdd.n1406 1.2505
R4406 avdd.n1405 avdd.n1404 1.2505
R4407 avdd.n1406 avdd.n1405 1.2505
R4408 avdd.n1205 avdd.n1203 1.2505
R4409 avdd.n1406 avdd.n1205 1.2505
R4410 avdd.n949 avdd.n932 1.16964
R4411 avdd.n947 avdd.n946 1.15136
R4412 avdd.n946 avdd.n945 1.15136
R4413 avdd.n945 avdd.n944 1.15136
R4414 avdd.n944 avdd.n943 1.15136
R4415 avdd.n943 avdd.n942 1.15136
R4416 avdd.n942 avdd.n941 1.15136
R4417 avdd.n939 avdd.n938 1.15136
R4418 avdd.n938 avdd.n937 1.15136
R4419 avdd.n937 avdd.n936 1.15136
R4420 avdd.n936 avdd.n935 1.15136
R4421 avdd.n935 avdd.n934 1.15136
R4422 avdd.n934 avdd.n933 1.15136
R4423 avdd.n933 avdd.n689 1.15136
R4424 avdd.n1018 avdd.n1015 1.14248
R4425 avdd.n1017 avdd.n1015 1.14248
R4426 avdd.n1016 avdd.n1014 1.14248
R4427 avdd.n1143 avdd.n1016 1.14248
R4428 avdd.n1264 avdd.n1261 1.14248
R4429 avdd.n1263 avdd.n1261 1.14248
R4430 avdd.n1262 avdd.n1260 1.14248
R4431 avdd.n1389 avdd.n1262 1.14248
R4432 avdd.n1650 avdd.n689 1.13628
R4433 avdd.n1486 avdd.n1454 1.12991
R4434 avdd.n941 avdd.n940 1.0824
R4435 avdd.n1063 avdd.n1062 1.05355
R4436 avdd.n1062 avdd.n952 1.05355
R4437 avdd.n1309 avdd.n1308 1.05355
R4438 avdd.n1308 avdd.n1198 1.05355
R4439 avdd.n1187 avdd.n1185 1.04347
R4440 avdd.n1055 avdd.n1053 1.04347
R4441 avdd.n995 avdd.n993 1.04347
R4442 avdd.n1089 avdd.n1065 1.04347
R4443 avdd.n1095 avdd.n1092 1.04347
R4444 avdd.n1433 avdd.n1431 1.04347
R4445 avdd.n1301 avdd.n1299 1.04347
R4446 avdd.n1241 avdd.n1239 1.04347
R4447 avdd.n1335 avdd.n1311 1.04347
R4448 avdd.n1341 avdd.n1338 1.04347
R4449 avdd.n1447 avdd.n951 1.03383
R4450 avdd.n1454 avdd.n1449 0.989805
R4451 avdd.n1493 avdd.n1449 0.989805
R4452 avdd.n672 avdd 0.983
R4453 avdd.n1469 avdd.n1468 0.954108
R4454 avdd.n1468 avdd.n1467 0.954108
R4455 avdd.n1541 avdd.n1539 0.907363
R4456 avdd.n1545 avdd.n1539 0.907363
R4457 avdd.n1542 avdd.n1540 0.907363
R4458 avdd.n1545 avdd.n1540 0.907363
R4459 avdd.n1639 avdd.n1606 0.90425
R4460 avdd.n1480 avdd.n1479 0.877277
R4461 avdd.n1479 avdd.n1478 0.877277
R4462 avdd avdd.n674 0.876125
R4463 avdd.n950 avdd.n949 0.83425
R4464 avdd.n1020 avdd.n1012 0.773938
R4465 avdd.n1266 avdd.n1258 0.773938
R4466 avdd.n125 avdd 0.755
R4467 avdd.n153 avdd 0.755
R4468 avdd.n181 avdd 0.755
R4469 avdd.n209 avdd 0.755
R4470 avdd.n237 avdd 0.755
R4471 avdd.n265 avdd 0.755
R4472 avdd.n293 avdd 0.755
R4473 avdd.n321 avdd 0.755
R4474 avdd.n461 avdd 0.755
R4475 avdd.n489 avdd 0.755
R4476 avdd.n517 avdd 0.755
R4477 avdd.n545 avdd 0.755
R4478 avdd.n573 avdd 0.755
R4479 avdd.n601 avdd 0.755
R4480 avdd.n629 avdd 0.755
R4481 avdd.n657 avdd 0.755
R4482 avdd.n1151 avdd.n1010 0.725109
R4483 avdd.n1397 avdd.n1256 0.725109
R4484 avdd.n1196 avdd.n1195 0.713391
R4485 avdd.n1193 avdd.n1191 0.713391
R4486 avdd.n1191 avdd.n1189 0.713391
R4487 avdd.n1189 avdd.n1187 0.713391
R4488 avdd.n1185 avdd.n1183 0.713391
R4489 avdd.n1183 avdd.n1181 0.713391
R4490 avdd.n1181 avdd.n1179 0.713391
R4491 avdd.n1179 avdd.n1177 0.713391
R4492 avdd.n1177 avdd.n1175 0.713391
R4493 avdd.n1175 avdd.n1173 0.713391
R4494 avdd.n1061 avdd.n1059 0.713391
R4495 avdd.n1059 avdd.n1057 0.713391
R4496 avdd.n1057 avdd.n1055 0.713391
R4497 avdd.n1053 avdd.n1051 0.713391
R4498 avdd.n1051 avdd.n1049 0.713391
R4499 avdd.n1049 avdd.n1047 0.713391
R4500 avdd.n1047 avdd.n1045 0.713391
R4501 avdd.n1045 avdd.n1043 0.713391
R4502 avdd.n1043 avdd.n982 0.713391
R4503 avdd.n989 avdd.n987 0.713391
R4504 avdd.n991 avdd.n989 0.713391
R4505 avdd.n993 avdd.n991 0.713391
R4506 avdd.n997 avdd.n995 0.713391
R4507 avdd.n999 avdd.n997 0.713391
R4508 avdd.n1001 avdd.n999 0.713391
R4509 avdd.n1003 avdd.n1001 0.713391
R4510 avdd.n1005 avdd.n1003 0.713391
R4511 avdd.n1007 avdd.n1005 0.713391
R4512 avdd.n1103 avdd.n1102 0.713391
R4513 avdd.n1102 avdd.n1099 0.713391
R4514 avdd.n1099 avdd.n1065 0.713391
R4515 avdd.n1089 avdd.n1088 0.713391
R4516 avdd.n1088 avdd.n1085 0.713391
R4517 avdd.n1085 avdd.n1067 0.713391
R4518 avdd.n1075 avdd.n1067 0.713391
R4519 avdd.n1075 avdd.n1074 0.713391
R4520 avdd.n1074 avdd.n1071 0.713391
R4521 avdd.n1106 avdd.n1064 0.713391
R4522 avdd.n1096 avdd.n1064 0.713391
R4523 avdd.n1096 avdd.n1095 0.713391
R4524 avdd.n1092 avdd.n1066 0.713391
R4525 avdd.n1082 avdd.n1066 0.713391
R4526 avdd.n1082 avdd.n1081 0.713391
R4527 avdd.n1081 avdd.n1078 0.713391
R4528 avdd.n1078 avdd.n1068 0.713391
R4529 avdd.n1068 avdd.n1025 0.713391
R4530 avdd.n1442 avdd.n1441 0.713391
R4531 avdd.n1439 avdd.n1437 0.713391
R4532 avdd.n1437 avdd.n1435 0.713391
R4533 avdd.n1435 avdd.n1433 0.713391
R4534 avdd.n1431 avdd.n1429 0.713391
R4535 avdd.n1429 avdd.n1427 0.713391
R4536 avdd.n1427 avdd.n1425 0.713391
R4537 avdd.n1425 avdd.n1423 0.713391
R4538 avdd.n1423 avdd.n1421 0.713391
R4539 avdd.n1421 avdd.n1419 0.713391
R4540 avdd.n1307 avdd.n1305 0.713391
R4541 avdd.n1305 avdd.n1303 0.713391
R4542 avdd.n1303 avdd.n1301 0.713391
R4543 avdd.n1299 avdd.n1297 0.713391
R4544 avdd.n1297 avdd.n1295 0.713391
R4545 avdd.n1295 avdd.n1293 0.713391
R4546 avdd.n1293 avdd.n1291 0.713391
R4547 avdd.n1291 avdd.n1289 0.713391
R4548 avdd.n1289 avdd.n1228 0.713391
R4549 avdd.n1235 avdd.n1233 0.713391
R4550 avdd.n1237 avdd.n1235 0.713391
R4551 avdd.n1239 avdd.n1237 0.713391
R4552 avdd.n1243 avdd.n1241 0.713391
R4553 avdd.n1245 avdd.n1243 0.713391
R4554 avdd.n1247 avdd.n1245 0.713391
R4555 avdd.n1249 avdd.n1247 0.713391
R4556 avdd.n1251 avdd.n1249 0.713391
R4557 avdd.n1253 avdd.n1251 0.713391
R4558 avdd.n1349 avdd.n1348 0.713391
R4559 avdd.n1348 avdd.n1345 0.713391
R4560 avdd.n1345 avdd.n1311 0.713391
R4561 avdd.n1335 avdd.n1334 0.713391
R4562 avdd.n1334 avdd.n1331 0.713391
R4563 avdd.n1331 avdd.n1313 0.713391
R4564 avdd.n1321 avdd.n1313 0.713391
R4565 avdd.n1321 avdd.n1320 0.713391
R4566 avdd.n1320 avdd.n1317 0.713391
R4567 avdd.n1352 avdd.n1310 0.713391
R4568 avdd.n1342 avdd.n1310 0.713391
R4569 avdd.n1342 avdd.n1341 0.713391
R4570 avdd.n1338 avdd.n1312 0.713391
R4571 avdd.n1328 avdd.n1312 0.713391
R4572 avdd.n1328 avdd.n1327 0.713391
R4573 avdd.n1327 avdd.n1324 0.713391
R4574 avdd.n1324 avdd.n1314 0.713391
R4575 avdd.n1314 avdd.n1271 0.713391
R4576 avdd.n1111 avdd.n1109 0.695812
R4577 avdd.n1113 avdd.n1111 0.695812
R4578 avdd.n1115 avdd.n1113 0.695812
R4579 avdd.n1117 avdd.n1115 0.695812
R4580 avdd.n1118 avdd.n1117 0.695812
R4581 avdd.n1357 avdd.n1355 0.695812
R4582 avdd.n1359 avdd.n1357 0.695812
R4583 avdd.n1361 avdd.n1359 0.695812
R4584 avdd.n1363 avdd.n1361 0.695812
R4585 avdd.n1364 avdd.n1363 0.695812
R4586 avdd.n77 avdd 0.664
R4587 avdd.n413 avdd 0.664
R4588 avdd.n1156 avdd.n1154 0.662609
R4589 avdd.n1402 avdd.n1400 0.662609
R4590 avdd.n1652 avdd.n1651 0.624875
R4591 avdd.n673 avdd 0.563625
R4592 avdd.n1457 avdd.n1456 0.56281
R4593 avdd.n1477 avdd.n1457 0.56281
R4594 avdd.n1463 avdd.n1448 0.559412
R4595 avdd.n1450 avdd.n1448 0.559412
R4596 avdd.n1640 avdd.n688 0.55425
R4597 avdd.n1576 avdd.n1575 0.545446
R4598 avdd.n1575 avdd.n1573 0.545446
R4599 avdd.n1573 avdd.n1571 0.545446
R4600 avdd.n1564 avdd.n1561 0.545446
R4601 avdd.n1557 avdd.n1556 0.545446
R4602 avdd.n1107 avdd.n1063 0.527027
R4603 avdd.n1194 avdd.n952 0.527027
R4604 avdd.n1353 avdd.n1309 0.527027
R4605 avdd.n1440 avdd.n1198 0.527027
R4606 avdd.n1173 avdd.n1171 0.477062
R4607 avdd.n1157 avdd.n982 0.477062
R4608 avdd.n1008 avdd.n1007 0.477062
R4609 avdd.n1071 avdd.n1024 0.477062
R4610 avdd.n1131 avdd.n1025 0.477062
R4611 avdd.n1419 avdd.n1417 0.477062
R4612 avdd.n1403 avdd.n1228 0.477062
R4613 avdd.n1254 avdd.n1253 0.477062
R4614 avdd.n1317 avdd.n1270 0.477062
R4615 avdd.n1377 avdd.n1271 0.477062
R4616 avdd.n1453 avdd.n1452 0.444145
R4617 avdd.n1452 avdd.n1451 0.444145
R4618 avdd.n1499 avdd.n1444 0.418878
R4619 avdd.n1502 avdd.n951 0.4145
R4620 avdd.n674 avdd.n673 0.407375
R4621 avdd.n1496 avdd.n1495 0.330857
R4622 avdd.n1495 avdd.n1494 0.330857
R4623 avdd.n1652 avdd 0.32398
R4624 avdd.n1171 avdd.n954 0.318859
R4625 avdd.n1157 avdd.n1156 0.318859
R4626 avdd.n1010 avdd.n1008 0.318859
R4627 avdd.n1135 avdd.n1024 0.318859
R4628 avdd.n1132 avdd.n1131 0.318859
R4629 avdd.n1417 avdd.n1200 0.318859
R4630 avdd.n1403 avdd.n1402 0.318859
R4631 avdd.n1256 avdd.n1254 0.318859
R4632 avdd.n1381 avdd.n1270 0.318859
R4633 avdd.n1378 avdd.n1377 0.318859
R4634 avdd.n1565 avdd.n1503 0.316162
R4635 avdd.n1531 avdd.n1529 0.291392
R4636 avdd.n1529 avdd.n1527 0.291392
R4637 avdd.n1551 avdd.n1550 0.284354
R4638 avdd.n1568 avdd.n1567 0.284354
R4639 avdd.n1651 avdd.n688 0.2805
R4640 avdd.n1565 avdd.n1564 0.273291
R4641 avdd.n1579 avdd.n1576 0.272973
R4642 avdd.n1561 avdd.n1557 0.272973
R4643 avdd.n1556 avdd.n1554 0.272973
R4644 avdd.n1109 avdd.n1108 0.262219
R4645 avdd.n1355 avdd.n1354 0.262219
R4646 avdd.n1502 avdd.n1501 0.2505
R4647 avdd avdd.n925 0.248811
R4648 avdd avdd.n914 0.248811
R4649 avdd.n717 avdd 0.248811
R4650 avdd avdd.n900 0.248811
R4651 avdd avdd.n889 0.248811
R4652 avdd.n737 avdd 0.248811
R4653 avdd avdd.n875 0.248811
R4654 avdd avdd.n864 0.248811
R4655 avdd.n757 avdd 0.248811
R4656 avdd avdd.n850 0.248811
R4657 avdd avdd.n839 0.248811
R4658 avdd.n777 avdd 0.248811
R4659 avdd avdd.n825 0.248811
R4660 avdd avdd.n814 0.248811
R4661 avdd.n797 avdd 0.248811
R4662 avdd.n1521 avdd.n1520 0.246297
R4663 avdd.n1500 avdd 0.242804
R4664 avdd.n1640 avdd.n1639 0.238625
R4665 avdd.n1571 avdd.n1503 0.229784
R4666 avdd.n1197 avdd.n1194 0.227878
R4667 avdd.n1443 avdd.n1440 0.227878
R4668 avdd.n1629 avdd.n1608 0.227329
R4669 avdd.n1636 avdd.n1635 0.227329
R4670 avdd.n1532 avdd.n1531 0.1885
R4671 avdd.n1471 avdd.n1470 0.1865
R4672 avdd.n1526 avdd.n1524 0.183736
R4673 avdd.n688 avdd.n687 0.175331
R4674 avdd.n1603 avdd.n1505 0.156108
R4675 avdd.n1148 avdd.n1147 0.152959
R4676 avdd.n1139 avdd.n1138 0.152959
R4677 avdd.n1394 avdd.n1393 0.152959
R4678 avdd.n1385 avdd.n1384 0.152959
R4679 avdd.n1489 avdd.n1488 0.152959
R4680 avdd.n1033 avdd.n1032 0.143577
R4681 avdd.n1279 avdd.n1278 0.143577
R4682 avdd.n1028 avdd.n1027 0.141409
R4683 avdd.n1274 avdd.n1273 0.141409
R4684 avdd.n1590 avdd.n1507 0.126176
R4685 avdd.n1595 avdd.n1506 0.126176
R4686 avdd.n1473 avdd.n1472 0.119731
R4687 avdd.n1611 avdd.n1607 0.113554
R4688 avdd.n1613 avdd.n1611 0.113554
R4689 avdd.n1615 avdd.n1613 0.113554
R4690 avdd.n1617 avdd.n1615 0.113554
R4691 avdd.n1619 avdd.n1617 0.113554
R4692 avdd.n1621 avdd.n1619 0.113554
R4693 avdd.n1623 avdd.n1621 0.113554
R4694 avdd.n1624 avdd.n1623 0.113554
R4695 avdd.n1524 avdd.n1523 0.113554
R4696 avdd.n1523 avdd.n1522 0.113554
R4697 avdd.n1566 avdd.n1552 0.0934054
R4698 avdd.n684 avdd.n676 0.0815811
R4699 avdd.n932 avdd.n696 0.0815811
R4700 avdd.n925 avdd.n701 0.0815811
R4701 avdd.n914 avdd.n708 0.0815811
R4702 avdd.n904 avdd.n717 0.0815811
R4703 avdd.n900 avdd.n720 0.0815811
R4704 avdd.n889 avdd.n728 0.0815811
R4705 avdd.n879 avdd.n737 0.0815811
R4706 avdd.n875 avdd.n740 0.0815811
R4707 avdd.n864 avdd.n748 0.0815811
R4708 avdd.n854 avdd.n757 0.0815811
R4709 avdd.n850 avdd.n760 0.0815811
R4710 avdd.n839 avdd.n768 0.0815811
R4711 avdd.n829 avdd.n777 0.0815811
R4712 avdd.n825 avdd.n780 0.0815811
R4713 avdd.n814 avdd.n788 0.0815811
R4714 avdd.n804 avdd.n797 0.0815811
R4715 avdd.n1642 avdd.n695 0.0793136
R4716 avdd.n940 avdd.n690 0.0793136
R4717 avdd.n1023 avdd.n1022 0.0766719
R4718 avdd.n1269 avdd.n1268 0.0766719
R4719 avdd.n940 avdd.n939 0.0694655
R4720 avdd.n1153 avdd.n957 0.0674065
R4721 avdd.n1399 avdd.n1203 0.0674065
R4722 avdd.n1162 avdd.n977 0.0669286
R4723 avdd.n1030 avdd.n964 0.0669286
R4724 avdd.n1408 avdd.n1223 0.0669286
R4725 avdd.n1276 avdd.n1210 0.0669286
R4726 avdd.n1022 avdd.n1019 0.0650833
R4727 avdd.n1013 avdd.n1012 0.0650833
R4728 avdd.n1268 avdd.n1265 0.0650833
R4729 avdd.n1259 avdd.n1258 0.0650833
R4730 avdd.n314 avdd.n312 0.0579519
R4731 avdd.n286 avdd.n284 0.0579519
R4732 avdd.n258 avdd.n256 0.0579519
R4733 avdd.n230 avdd.n228 0.0579519
R4734 avdd.n202 avdd.n200 0.0579519
R4735 avdd.n174 avdd.n172 0.0579519
R4736 avdd.n146 avdd.n144 0.0579519
R4737 avdd.n118 avdd.n116 0.0579519
R4738 avdd.n87 avdd.n83 0.0579519
R4739 avdd.n650 avdd.n648 0.0579519
R4740 avdd.n622 avdd.n620 0.0579519
R4741 avdd.n594 avdd.n592 0.0579519
R4742 avdd.n566 avdd.n564 0.0579519
R4743 avdd.n538 avdd.n536 0.0579519
R4744 avdd.n510 avdd.n508 0.0579519
R4745 avdd.n482 avdd.n480 0.0579519
R4746 avdd.n454 avdd.n452 0.0579519
R4747 avdd.n423 avdd.n419 0.0579519
R4748 avdd.n685 avdd.n675 0.0553986
R4749 avdd.n928 avdd.n700 0.0553986
R4750 avdd.n917 avdd.n707 0.0553986
R4751 avdd.n714 avdd.n713 0.0553986
R4752 avdd.n903 avdd.n719 0.0553986
R4753 avdd.n892 avdd.n727 0.0553986
R4754 avdd.n734 avdd.n733 0.0553986
R4755 avdd.n878 avdd.n739 0.0553986
R4756 avdd.n867 avdd.n747 0.0553986
R4757 avdd.n754 avdd.n753 0.0553986
R4758 avdd.n853 avdd.n759 0.0553986
R4759 avdd.n842 avdd.n767 0.0553986
R4760 avdd.n774 avdd.n773 0.0553986
R4761 avdd.n828 avdd.n779 0.0553986
R4762 avdd.n817 avdd.n787 0.0553986
R4763 avdd.n794 avdd.n793 0.0553986
R4764 avdd.n803 avdd.n800 0.0553986
R4765 avdd.n1487 avdd.n1486 0.0527472
R4766 avdd.n1485 avdd.n1484 0.0510435
R4767 avdd.n1466 avdd.n1462 0.0507703
R4768 avdd.n1543 avdd.n1541 0.0489375
R4769 avdd.n1569 avdd.n1542 0.0489375
R4770 avdd.n1482 avdd.n1481 0.0467687
R4771 avdd avdd.n1652 0.04675
R4772 avdd.n1527 avdd.n1526 0.0436892
R4773 avdd.n1638 avdd.n1607 0.0430541
R4774 avdd.n1532 avdd.n1521 0.0430541
R4775 avdd.n676 avdd 0.0410405
R4776 avdd avdd.n89 0.04
R4777 avdd avdd.n123 0.04
R4778 avdd avdd.n151 0.04
R4779 avdd avdd.n179 0.04
R4780 avdd avdd.n207 0.04
R4781 avdd avdd.n235 0.04
R4782 avdd avdd.n263 0.04
R4783 avdd avdd.n291 0.04
R4784 avdd avdd.n319 0.04
R4785 avdd avdd.n425 0.04
R4786 avdd avdd.n459 0.04
R4787 avdd avdd.n487 0.04
R4788 avdd avdd.n515 0.04
R4789 avdd avdd.n543 0.04
R4790 avdd avdd.n571 0.04
R4791 avdd avdd.n599 0.04
R4792 avdd avdd.n627 0.04
R4793 avdd avdd.n655 0.04
R4794 avdd.n1445 avdd.n951 0.0375
R4795 avdd avdd.n85 0.0365
R4796 avdd avdd.n114 0.0365
R4797 avdd avdd.n142 0.0365
R4798 avdd avdd.n170 0.0365
R4799 avdd avdd.n198 0.0365
R4800 avdd avdd.n226 0.0365
R4801 avdd avdd.n254 0.0365
R4802 avdd avdd.n282 0.0365
R4803 avdd avdd.n310 0.0365
R4804 avdd avdd.n421 0.0365
R4805 avdd avdd.n450 0.0365
R4806 avdd avdd.n478 0.0365
R4807 avdd avdd.n506 0.0365
R4808 avdd avdd.n534 0.0365
R4809 avdd avdd.n562 0.0365
R4810 avdd avdd.n590 0.0365
R4811 avdd avdd.n618 0.0365
R4812 avdd avdd.n646 0.0365
R4813 avdd.n927 avdd 0.0351284
R4814 avdd.n916 avdd 0.0351284
R4815 avdd avdd.n716 0.0351284
R4816 avdd.n901 avdd 0.0351284
R4817 avdd.n891 avdd 0.0351284
R4818 avdd avdd.n736 0.0351284
R4819 avdd.n876 avdd 0.0351284
R4820 avdd.n866 avdd 0.0351284
R4821 avdd avdd.n756 0.0351284
R4822 avdd.n851 avdd 0.0351284
R4823 avdd.n841 avdd 0.0351284
R4824 avdd avdd.n776 0.0351284
R4825 avdd.n826 avdd 0.0351284
R4826 avdd.n816 avdd 0.0351284
R4827 avdd avdd.n796 0.0351284
R4828 avdd.n801 avdd 0.0351284
R4829 avdd.n74 avdd 0.0335784
R4830 avdd.n410 avdd 0.0335784
R4831 avdd.n105 avdd 0.032
R4832 avdd.n133 avdd 0.032
R4833 avdd.n161 avdd 0.032
R4834 avdd.n189 avdd 0.032
R4835 avdd.n217 avdd 0.032
R4836 avdd.n245 avdd 0.032
R4837 avdd.n273 avdd 0.032
R4838 avdd.n301 avdd 0.032
R4839 avdd.n329 avdd 0.032
R4840 avdd.n441 avdd 0.032
R4841 avdd.n469 avdd 0.032
R4842 avdd.n497 avdd 0.032
R4843 avdd.n525 avdd 0.032
R4844 avdd.n553 avdd 0.032
R4845 avdd.n581 avdd 0.032
R4846 avdd.n609 avdd 0.032
R4847 avdd.n637 avdd 0.032
R4848 avdd.n665 avdd 0.032
R4849 avdd.n1461 avdd.n1455 0.0301178
R4850 avdd.n1465 avdd.n1464 0.0300238
R4851 avdd.n1522 avdd.n1505 0.0287635
R4852 avdd.n1498 avdd.n1497 0.0283443
R4853 avdd.n80 avdd 0.028
R4854 avdd.n416 avdd 0.028
R4855 avdd.n685 avdd.n684 0.0266824
R4856 avdd.n700 avdd.n696 0.0266824
R4857 avdd.n707 avdd.n701 0.0266824
R4858 avdd.n714 avdd.n708 0.0266824
R4859 avdd.n904 avdd.n903 0.0266824
R4860 avdd.n727 avdd.n720 0.0266824
R4861 avdd.n734 avdd.n728 0.0266824
R4862 avdd.n879 avdd.n878 0.0266824
R4863 avdd.n747 avdd.n740 0.0266824
R4864 avdd.n754 avdd.n748 0.0266824
R4865 avdd.n854 avdd.n853 0.0266824
R4866 avdd.n767 avdd.n760 0.0266824
R4867 avdd.n774 avdd.n768 0.0266824
R4868 avdd.n829 avdd.n828 0.0266824
R4869 avdd.n787 avdd.n780 0.0266824
R4870 avdd.n794 avdd.n788 0.0266824
R4871 avdd.n804 avdd.n803 0.0266824
R4872 avdd.n90 avdd 0.0245
R4873 avdd.n84 avdd 0.0245
R4874 avdd avdd.n124 0.0245
R4875 avdd.n120 avdd 0.0245
R4876 avdd avdd.n152 0.0245
R4877 avdd.n148 avdd 0.0245
R4878 avdd avdd.n180 0.0245
R4879 avdd.n176 avdd 0.0245
R4880 avdd avdd.n208 0.0245
R4881 avdd.n204 avdd 0.0245
R4882 avdd avdd.n236 0.0245
R4883 avdd.n232 avdd 0.0245
R4884 avdd avdd.n264 0.0245
R4885 avdd.n260 avdd 0.0245
R4886 avdd avdd.n292 0.0245
R4887 avdd.n288 avdd 0.0245
R4888 avdd avdd.n320 0.0245
R4889 avdd.n316 avdd 0.0245
R4890 avdd.n420 avdd 0.0245
R4891 avdd avdd.n460 0.0245
R4892 avdd.n456 avdd 0.0245
R4893 avdd avdd.n488 0.0245
R4894 avdd.n484 avdd 0.0245
R4895 avdd avdd.n516 0.0245
R4896 avdd.n512 avdd 0.0245
R4897 avdd avdd.n544 0.0245
R4898 avdd.n540 avdd 0.0245
R4899 avdd avdd.n572 0.0245
R4900 avdd.n568 avdd 0.0245
R4901 avdd avdd.n600 0.0245
R4902 avdd.n596 avdd 0.0245
R4903 avdd avdd.n628 0.0245
R4904 avdd.n624 avdd 0.0245
R4905 avdd avdd.n656 0.0245
R4906 avdd.n652 avdd 0.0245
R4907 avdd.n1483 avdd.n1453 0.0240443
R4908 avdd.n426 avdd 0.024
R4909 avdd avdd.n74 0.0163924
R4910 avdd avdd.n410 0.0163924
R4911 avdd avdd.n1197 0.01225
R4912 avdd avdd.n1443 0.01225
R4913 avdd avdd.n64 0.012
R4914 avdd avdd.n56 0.012
R4915 avdd avdd.n48 0.012
R4916 avdd avdd.n40 0.012
R4917 avdd avdd.n32 0.012
R4918 avdd avdd.n24 0.012
R4919 avdd avdd.n16 0.012
R4920 avdd avdd.n8 0.012
R4921 avdd avdd.n0 0.012
R4922 avdd avdd.n400 0.012
R4923 avdd avdd.n392 0.012
R4924 avdd avdd.n384 0.012
R4925 avdd avdd.n376 0.012
R4926 avdd avdd.n368 0.012
R4927 avdd avdd.n360 0.012
R4928 avdd avdd.n352 0.012
R4929 avdd avdd.n344 0.012
R4930 avdd avdd.n336 0.012
R4931 avdd avdd.n77 0.009
R4932 avdd.n78 avdd 0.009
R4933 avdd.n90 avdd 0.009
R4934 avdd.n89 avdd 0.009
R4935 avdd.n88 avdd 0.009
R4936 avdd.n85 avdd 0.009
R4937 avdd.n109 avdd 0.009
R4938 avdd.n109 avdd 0.009
R4939 avdd.n108 avdd 0.009
R4940 avdd.n125 avdd 0.009
R4941 avdd.n124 avdd 0.009
R4942 avdd.n123 avdd 0.009
R4943 avdd.n117 avdd 0.009
R4944 avdd.n114 avdd 0.009
R4945 avdd.n137 avdd 0.009
R4946 avdd.n137 avdd 0.009
R4947 avdd.n136 avdd 0.009
R4948 avdd.n153 avdd 0.009
R4949 avdd.n152 avdd 0.009
R4950 avdd.n151 avdd 0.009
R4951 avdd.n145 avdd 0.009
R4952 avdd.n142 avdd 0.009
R4953 avdd.n165 avdd 0.009
R4954 avdd.n165 avdd 0.009
R4955 avdd.n164 avdd 0.009
R4956 avdd.n181 avdd 0.009
R4957 avdd.n180 avdd 0.009
R4958 avdd.n179 avdd 0.009
R4959 avdd.n173 avdd 0.009
R4960 avdd.n170 avdd 0.009
R4961 avdd.n193 avdd 0.009
R4962 avdd.n193 avdd 0.009
R4963 avdd.n192 avdd 0.009
R4964 avdd.n209 avdd 0.009
R4965 avdd.n208 avdd 0.009
R4966 avdd.n207 avdd 0.009
R4967 avdd.n201 avdd 0.009
R4968 avdd.n198 avdd 0.009
R4969 avdd.n221 avdd 0.009
R4970 avdd.n221 avdd 0.009
R4971 avdd.n220 avdd 0.009
R4972 avdd.n237 avdd 0.009
R4973 avdd.n236 avdd 0.009
R4974 avdd.n235 avdd 0.009
R4975 avdd.n229 avdd 0.009
R4976 avdd.n226 avdd 0.009
R4977 avdd.n249 avdd 0.009
R4978 avdd.n249 avdd 0.009
R4979 avdd.n248 avdd 0.009
R4980 avdd.n265 avdd 0.009
R4981 avdd.n264 avdd 0.009
R4982 avdd.n263 avdd 0.009
R4983 avdd.n257 avdd 0.009
R4984 avdd.n254 avdd 0.009
R4985 avdd.n277 avdd 0.009
R4986 avdd.n277 avdd 0.009
R4987 avdd.n276 avdd 0.009
R4988 avdd.n293 avdd 0.009
R4989 avdd.n292 avdd 0.009
R4990 avdd.n291 avdd 0.009
R4991 avdd.n285 avdd 0.009
R4992 avdd.n282 avdd 0.009
R4993 avdd.n305 avdd 0.009
R4994 avdd.n305 avdd 0.009
R4995 avdd.n304 avdd 0.009
R4996 avdd.n321 avdd 0.009
R4997 avdd.n320 avdd 0.009
R4998 avdd.n319 avdd 0.009
R4999 avdd.n313 avdd 0.009
R5000 avdd.n310 avdd 0.009
R5001 avdd.n333 avdd 0.009
R5002 avdd.n333 avdd 0.009
R5003 avdd.n332 avdd 0.009
R5004 avdd avdd.n413 0.009
R5005 avdd.n414 avdd 0.009
R5006 avdd.n426 avdd 0.009
R5007 avdd.n425 avdd 0.009
R5008 avdd.n424 avdd 0.009
R5009 avdd.n421 avdd 0.009
R5010 avdd.n445 avdd 0.009
R5011 avdd.n445 avdd 0.009
R5012 avdd.n444 avdd 0.009
R5013 avdd.n461 avdd 0.009
R5014 avdd.n460 avdd 0.009
R5015 avdd.n459 avdd 0.009
R5016 avdd.n453 avdd 0.009
R5017 avdd.n450 avdd 0.009
R5018 avdd.n473 avdd 0.009
R5019 avdd.n473 avdd 0.009
R5020 avdd.n472 avdd 0.009
R5021 avdd.n489 avdd 0.009
R5022 avdd.n488 avdd 0.009
R5023 avdd.n487 avdd 0.009
R5024 avdd.n481 avdd 0.009
R5025 avdd.n478 avdd 0.009
R5026 avdd.n501 avdd 0.009
R5027 avdd.n501 avdd 0.009
R5028 avdd.n500 avdd 0.009
R5029 avdd.n517 avdd 0.009
R5030 avdd.n516 avdd 0.009
R5031 avdd.n515 avdd 0.009
R5032 avdd.n509 avdd 0.009
R5033 avdd.n506 avdd 0.009
R5034 avdd.n529 avdd 0.009
R5035 avdd.n529 avdd 0.009
R5036 avdd.n528 avdd 0.009
R5037 avdd.n545 avdd 0.009
R5038 avdd.n544 avdd 0.009
R5039 avdd.n543 avdd 0.009
R5040 avdd.n537 avdd 0.009
R5041 avdd.n534 avdd 0.009
R5042 avdd.n557 avdd 0.009
R5043 avdd.n557 avdd 0.009
R5044 avdd.n556 avdd 0.009
R5045 avdd.n573 avdd 0.009
R5046 avdd.n572 avdd 0.009
R5047 avdd.n571 avdd 0.009
R5048 avdd.n565 avdd 0.009
R5049 avdd.n562 avdd 0.009
R5050 avdd.n585 avdd 0.009
R5051 avdd.n585 avdd 0.009
R5052 avdd.n584 avdd 0.009
R5053 avdd.n601 avdd 0.009
R5054 avdd.n600 avdd 0.009
R5055 avdd.n599 avdd 0.009
R5056 avdd.n593 avdd 0.009
R5057 avdd.n590 avdd 0.009
R5058 avdd.n613 avdd 0.009
R5059 avdd.n613 avdd 0.009
R5060 avdd.n612 avdd 0.009
R5061 avdd.n629 avdd 0.009
R5062 avdd.n628 avdd 0.009
R5063 avdd.n627 avdd 0.009
R5064 avdd.n621 avdd 0.009
R5065 avdd.n618 avdd 0.009
R5066 avdd.n641 avdd 0.009
R5067 avdd.n641 avdd 0.009
R5068 avdd.n640 avdd 0.009
R5069 avdd.n657 avdd 0.009
R5070 avdd.n656 avdd 0.009
R5071 avdd.n655 avdd 0.009
R5072 avdd.n649 avdd 0.009
R5073 avdd.n646 avdd 0.009
R5074 avdd.n669 avdd 0.009
R5075 avdd.n669 avdd 0.009
R5076 avdd.n668 avdd 0.009
R5077 avdd avdd.n81 0.0085
R5078 avdd.n105 avdd.n104 0.0085
R5079 avdd.n133 avdd.n132 0.0085
R5080 avdd.n161 avdd.n160 0.0085
R5081 avdd.n189 avdd.n188 0.0085
R5082 avdd.n217 avdd.n216 0.0085
R5083 avdd.n245 avdd.n244 0.0085
R5084 avdd.n273 avdd.n272 0.0085
R5085 avdd.n301 avdd.n300 0.0085
R5086 avdd.n329 avdd.n328 0.0085
R5087 avdd avdd.n417 0.0085
R5088 avdd.n441 avdd.n440 0.0085
R5089 avdd.n469 avdd.n468 0.0085
R5090 avdd.n497 avdd.n496 0.0085
R5091 avdd.n525 avdd.n524 0.0085
R5092 avdd.n553 avdd.n552 0.0085
R5093 avdd.n581 avdd.n580 0.0085
R5094 avdd.n609 avdd.n608 0.0085
R5095 avdd.n637 avdd.n636 0.0085
R5096 avdd.n665 avdd.n664 0.0085
R5097 avdd avdd.n88 0.0075
R5098 avdd.n117 avdd 0.0075
R5099 avdd.n145 avdd 0.0075
R5100 avdd.n173 avdd 0.0075
R5101 avdd.n201 avdd 0.0075
R5102 avdd.n229 avdd 0.0075
R5103 avdd.n257 avdd 0.0075
R5104 avdd.n285 avdd 0.0075
R5105 avdd.n313 avdd 0.0075
R5106 avdd avdd.n424 0.0075
R5107 avdd.n453 avdd 0.0075
R5108 avdd.n481 avdd 0.0075
R5109 avdd.n509 avdd 0.0075
R5110 avdd.n537 avdd 0.0075
R5111 avdd.n565 avdd 0.0075
R5112 avdd.n593 avdd 0.0075
R5113 avdd.n621 avdd 0.0075
R5114 avdd.n649 avdd 0.0075
R5115 avdd.n687 avdd.n675 0.00641216
R5116 avdd.n928 avdd.n927 0.00641216
R5117 avdd.n917 avdd.n916 0.00641216
R5118 avdd.n716 avdd.n713 0.00641216
R5119 avdd.n901 avdd.n719 0.00641216
R5120 avdd.n892 avdd.n891 0.00641216
R5121 avdd.n736 avdd.n733 0.00641216
R5122 avdd.n876 avdd.n739 0.00641216
R5123 avdd.n867 avdd.n866 0.00641216
R5124 avdd.n756 avdd.n753 0.00641216
R5125 avdd.n851 avdd.n759 0.00641216
R5126 avdd.n842 avdd.n841 0.00641216
R5127 avdd.n776 avdd.n773 0.00641216
R5128 avdd.n826 avdd.n779 0.00641216
R5129 avdd.n817 avdd.n816 0.00641216
R5130 avdd.n796 avdd.n793 0.00641216
R5131 avdd.n801 avdd.n800 0.00641216
R5132 avdd.n86 avdd 0.0055
R5133 avdd.n111 avdd.n64 0.0055
R5134 avdd.n119 avdd 0.0055
R5135 avdd.n139 avdd.n56 0.0055
R5136 avdd.n147 avdd 0.0055
R5137 avdd.n167 avdd.n48 0.0055
R5138 avdd.n175 avdd 0.0055
R5139 avdd.n195 avdd.n40 0.0055
R5140 avdd.n203 avdd 0.0055
R5141 avdd.n223 avdd.n32 0.0055
R5142 avdd.n231 avdd 0.0055
R5143 avdd.n251 avdd.n24 0.0055
R5144 avdd.n259 avdd 0.0055
R5145 avdd.n279 avdd.n16 0.0055
R5146 avdd.n287 avdd 0.0055
R5147 avdd.n307 avdd.n8 0.0055
R5148 avdd.n315 avdd 0.0055
R5149 avdd.n335 avdd.n0 0.0055
R5150 avdd.n422 avdd 0.0055
R5151 avdd.n447 avdd.n400 0.0055
R5152 avdd.n455 avdd 0.0055
R5153 avdd.n475 avdd.n392 0.0055
R5154 avdd.n483 avdd 0.0055
R5155 avdd.n503 avdd.n384 0.0055
R5156 avdd.n511 avdd 0.0055
R5157 avdd.n531 avdd.n376 0.0055
R5158 avdd.n539 avdd 0.0055
R5159 avdd.n559 avdd.n368 0.0055
R5160 avdd.n567 avdd 0.0055
R5161 avdd.n587 avdd.n360 0.0055
R5162 avdd.n595 avdd 0.0055
R5163 avdd.n615 avdd.n352 0.0055
R5164 avdd.n623 avdd 0.0055
R5165 avdd.n643 avdd.n344 0.0055
R5166 avdd.n651 avdd 0.0055
R5167 avdd.n671 avdd.n336 0.0055
R5168 avdd.n86 avdd.n84 0.004
R5169 avdd avdd.n111 0.004
R5170 avdd.n120 avdd.n119 0.004
R5171 avdd avdd.n139 0.004
R5172 avdd.n148 avdd.n147 0.004
R5173 avdd avdd.n167 0.004
R5174 avdd.n176 avdd.n175 0.004
R5175 avdd avdd.n195 0.004
R5176 avdd.n204 avdd.n203 0.004
R5177 avdd avdd.n223 0.004
R5178 avdd.n232 avdd.n231 0.004
R5179 avdd avdd.n251 0.004
R5180 avdd.n260 avdd.n259 0.004
R5181 avdd avdd.n279 0.004
R5182 avdd.n288 avdd.n287 0.004
R5183 avdd avdd.n307 0.004
R5184 avdd.n316 avdd.n315 0.004
R5185 avdd avdd.n335 0.004
R5186 avdd.n422 avdd.n420 0.004
R5187 avdd avdd.n447 0.004
R5188 avdd.n456 avdd.n455 0.004
R5189 avdd avdd.n475 0.004
R5190 avdd.n484 avdd.n483 0.004
R5191 avdd avdd.n503 0.004
R5192 avdd.n512 avdd.n511 0.004
R5193 avdd avdd.n531 0.004
R5194 avdd.n540 avdd.n539 0.004
R5195 avdd avdd.n559 0.004
R5196 avdd.n568 avdd.n567 0.004
R5197 avdd avdd.n587 0.004
R5198 avdd.n596 avdd.n595 0.004
R5199 avdd avdd.n615 0.004
R5200 avdd.n624 avdd.n623 0.004
R5201 avdd avdd.n643 0.004
R5202 avdd.n652 avdd.n651 0.004
R5203 avdd avdd.n671 0.004
R5204 avdd.n78 avdd 0.0035
R5205 avdd.n414 avdd 0.0035
R5206 avdd avdd.n108 0.003
R5207 avdd avdd.n136 0.003
R5208 avdd avdd.n164 0.003
R5209 avdd avdd.n192 0.003
R5210 avdd avdd.n220 0.003
R5211 avdd avdd.n248 0.003
R5212 avdd avdd.n276 0.003
R5213 avdd avdd.n304 0.003
R5214 avdd avdd.n332 0.003
R5215 avdd avdd.n444 0.003
R5216 avdd avdd.n472 0.003
R5217 avdd avdd.n500 0.003
R5218 avdd avdd.n528 0.003
R5219 avdd avdd.n556 0.003
R5220 avdd avdd.n584 0.003
R5221 avdd avdd.n612 0.003
R5222 avdd avdd.n640 0.003
R5223 avdd avdd.n668 0.003
R5224 avdd.n81 avdd.n80 0.001
R5225 avdd.n104 avdd 0.001
R5226 avdd.n132 avdd 0.001
R5227 avdd.n160 avdd 0.001
R5228 avdd.n188 avdd 0.001
R5229 avdd.n216 avdd 0.001
R5230 avdd.n244 avdd 0.001
R5231 avdd.n272 avdd 0.001
R5232 avdd.n300 avdd 0.001
R5233 avdd.n328 avdd 0.001
R5234 avdd.n417 avdd.n416 0.001
R5235 avdd.n440 avdd 0.001
R5236 avdd.n468 avdd 0.001
R5237 avdd.n496 avdd 0.001
R5238 avdd.n524 avdd 0.001
R5239 avdd.n552 avdd 0.001
R5240 avdd.n580 avdd 0.001
R5241 avdd.n608 avdd 0.001
R5242 avdd.n636 avdd 0.001
R5243 avdd.n664 avdd 0.001
R5244 vunder.n2 vunder.n0 243.458
R5245 vunder.n2 vunder.n1 205.059
R5246 vunder.n4 vunder.n3 205.059
R5247 vunder.n6 vunder.n5 205.059
R5248 vunder.n8 vunder.n7 205.059
R5249 vunder.n10 vunder.n9 205.059
R5250 vunder.n12 vunder.n11 205.059
R5251 vunder.n14 vunder.n13 205.059
R5252 vunder.n17 vunder.n15 133.534
R5253 vunder.n17 vunder.n16 99.1759
R5254 vunder.n19 vunder.n18 99.1759
R5255 vunder.n21 vunder.n20 99.1759
R5256 vunder.n23 vunder.n22 99.1759
R5257 vunder.n25 vunder.n24 99.1759
R5258 vunder.n27 vunder.n26 99.1759
R5259 vunder vunder.n28 97.4305
R5260 vunder.n4 vunder.n2 38.4005
R5261 vunder.n6 vunder.n4 38.4005
R5262 vunder.n8 vunder.n6 38.4005
R5263 vunder.n10 vunder.n8 38.4005
R5264 vunder.n12 vunder.n10 38.4005
R5265 vunder.n14 vunder.n12 38.4005
R5266 vunder.n19 vunder.n17 34.3584
R5267 vunder.n21 vunder.n19 34.3584
R5268 vunder.n23 vunder.n21 34.3584
R5269 vunder.n25 vunder.n23 34.3584
R5270 vunder.n27 vunder.n25 34.3584
R5271 vunder.n29 vunder.n27 34.3584
R5272 vunder.n13 vunder.t1 26.5955
R5273 vunder.n13 vunder.t13 26.5955
R5274 vunder.n0 vunder.t2 26.5955
R5275 vunder.n0 vunder.t4 26.5955
R5276 vunder.n1 vunder.t8 26.5955
R5277 vunder.n1 vunder.t15 26.5955
R5278 vunder.n3 vunder.t12 26.5955
R5279 vunder.n3 vunder.t14 26.5955
R5280 vunder.n5 vunder.t11 26.5955
R5281 vunder.n5 vunder.t6 26.5955
R5282 vunder.n7 vunder.t0 26.5955
R5283 vunder.n7 vunder.t5 26.5955
R5284 vunder.n9 vunder.t10 26.5955
R5285 vunder.n9 vunder.t3 26.5955
R5286 vunder.n11 vunder.t9 26.5955
R5287 vunder.n11 vunder.t7 26.5955
R5288 vunder.n28 vunder.t29 24.9236
R5289 vunder.n28 vunder.t18 24.9236
R5290 vunder.n15 vunder.t27 24.9236
R5291 vunder.n15 vunder.t22 24.9236
R5292 vunder.n16 vunder.t26 24.9236
R5293 vunder.n16 vunder.t20 24.9236
R5294 vunder.n18 vunder.t17 24.9236
R5295 vunder.n18 vunder.t19 24.9236
R5296 vunder.n20 vunder.t16 24.9236
R5297 vunder.n20 vunder.t24 24.9236
R5298 vunder.n22 vunder.t28 24.9236
R5299 vunder.n22 vunder.t23 24.9236
R5300 vunder.n24 vunder.t31 24.9236
R5301 vunder.n24 vunder.t21 24.9236
R5302 vunder.n26 vunder.t30 24.9236
R5303 vunder.n26 vunder.t25 24.9236
R5304 vunder vunder.n14 18.4247
R5305 vunder.n30 vunder.n29 8.33989
R5306 vunder.n30 vunder 4.78765
R5307 vunder vunder.n30 3.10353
R5308 vunder.n29 vunder 1.74595
R5309 dvdd.n470 dvdd.n468 51406.3
R5310 dvdd.n472 dvdd.n468 51406.3
R5311 dvdd.n472 dvdd.n471 51406.3
R5312 dvdd.n471 dvdd.n470 51406.3
R5313 dvdd.n469 dvdd.n467 25491.9
R5314 dvdd.n473 dvdd.n467 25491.9
R5315 dvdd.n473 dvdd.n466 25491.9
R5316 dvdd.n469 dvdd.n466 25491.9
R5317 dvdd.n273 dvdd.n271 21292
R5318 dvdd.n274 dvdd.n273 21288.6
R5319 dvdd.n275 dvdd.n271 21288.6
R5320 dvdd.n275 dvdd.n274 21285.3
R5321 dvdd.n272 dvdd.n269 10790.3
R5322 dvdd.n272 dvdd.n270 10788.6
R5323 dvdd.n276 dvdd.n269 10788.6
R5324 dvdd.n276 dvdd.n270 10787
R5325 dvdd.n502 dvdd.n499 8474.12
R5326 dvdd.n504 dvdd.n499 8474.12
R5327 dvdd.n502 dvdd.n501 8470.59
R5328 dvdd.n504 dvdd.n501 8470.59
R5329 dvdd.n465 dvdd.n464 5925.65
R5330 dvdd.n475 dvdd.n465 5925.65
R5331 dvdd.n474 dvdd.n464 5925.65
R5332 dvdd.n475 dvdd.n474 5925.65
R5333 dvdd.n204 dvdd.n203 4782.35
R5334 dvdd.n205 dvdd.n203 4782.35
R5335 dvdd.n204 dvdd.n188 4782.35
R5336 dvdd.n205 dvdd.n188 4782.35
R5337 dvdd.n278 dvdd.n268 2512.56
R5338 dvdd.n268 dvdd.n267 2512.19
R5339 dvdd.n278 dvdd.n277 2512.19
R5340 dvdd.n277 dvdd.n267 2511.81
R5341 dvdd.n507 dvdd.n498 903.907
R5342 dvdd.n505 dvdd.n500 903.529
R5343 dvdd.n500 dvdd.n498 903.529
R5344 dvdd.n258 dvdd.t109 871.962
R5345 dvdd.n119 dvdd.t180 871.962
R5346 dvdd.n175 dvdd.t73 871.962
R5347 dvdd.n342 dvdd.t49 871.962
R5348 dvdd.n288 dvdd.t231 871.962
R5349 dvdd.n506 dvdd.n505 857.977
R5350 dvdd.n206 dvdd.n202 510.118
R5351 dvdd.n207 dvdd.n206 510.118
R5352 dvdd.n207 dvdd.n187 510.118
R5353 dvdd.n202 dvdd.n187 510.118
R5354 dvdd.t42 dvdd.n204 369.05
R5355 dvdd.n205 dvdd.t82 369.05
R5356 dvdd.n488 dvdd.t124 360.925
R5357 dvdd.n486 dvdd.t114 360.795
R5358 dvdd dvdd.t230 350
R5359 dvdd dvdd.t48 350
R5360 dvdd.n300 dvdd.t249 349.238
R5361 dvdd.n225 dvdd.t15 348.805
R5362 dvdd.n86 dvdd.t166 348.755
R5363 dvdd.n142 dvdd.t311 348.755
R5364 dvdd dvdd.t179 341.488
R5365 dvdd dvdd.t72 341.488
R5366 dvdd dvdd.t108 336.933
R5367 dvdd.n263 dvdd.n212 320.976
R5368 dvdd.n252 dvdd.n216 320.976
R5369 dvdd.n218 dvdd.n217 320.976
R5370 dvdd.n244 dvdd.n220 320.976
R5371 dvdd.n238 dvdd.n237 320.976
R5372 dvdd.n235 dvdd.n223 320.976
R5373 dvdd.n229 dvdd.n228 320.976
R5374 dvdd.n227 dvdd.n226 320.976
R5375 dvdd.n124 dvdd.n73 320.976
R5376 dvdd.n113 dvdd.n77 320.976
R5377 dvdd.n79 dvdd.n78 320.976
R5378 dvdd.n105 dvdd.n81 320.976
R5379 dvdd.n99 dvdd.n98 320.976
R5380 dvdd.n96 dvdd.n84 320.976
R5381 dvdd.n90 dvdd.n89 320.976
R5382 dvdd.n88 dvdd.n87 320.976
R5383 dvdd.n180 dvdd.n129 320.976
R5384 dvdd.n169 dvdd.n133 320.976
R5385 dvdd.n135 dvdd.n134 320.976
R5386 dvdd.n161 dvdd.n137 320.976
R5387 dvdd.n155 dvdd.n154 320.976
R5388 dvdd.n152 dvdd.n140 320.976
R5389 dvdd.n146 dvdd.n145 320.976
R5390 dvdd.n144 dvdd.n143 320.976
R5391 dvdd.n337 dvdd.n287 320.976
R5392 dvdd.n347 dvdd.n283 320.976
R5393 dvdd.n327 dvdd.n291 320.976
R5394 dvdd.n293 dvdd.n292 320.976
R5395 dvdd.n319 dvdd.n295 320.976
R5396 dvdd.n313 dvdd.n312 320.976
R5397 dvdd.n310 dvdd.n298 320.976
R5398 dvdd.n304 dvdd.n303 320.976
R5399 dvdd.n302 dvdd.n301 320.976
R5400 dvdd.n458 dvdd.n352 307.762
R5401 dvdd.n454 dvdd.n359 307.762
R5402 dvdd.n450 dvdd.n366 307.762
R5403 dvdd.n446 dvdd.n373 307.762
R5404 dvdd.n442 dvdd.n380 307.762
R5405 dvdd.n438 dvdd.n387 307.762
R5406 dvdd.n434 dvdd.n394 307.762
R5407 dvdd.n430 dvdd.n401 307.762
R5408 dvdd.n426 dvdd.n408 307.762
R5409 dvdd.n517 dvdd.n71 307.762
R5410 dvdd.n521 dvdd.n64 307.762
R5411 dvdd.n525 dvdd.n57 307.762
R5412 dvdd.n529 dvdd.n50 307.762
R5413 dvdd.n533 dvdd.n43 307.762
R5414 dvdd.n537 dvdd.n36 307.762
R5415 dvdd.n541 dvdd.n29 307.762
R5416 dvdd.n545 dvdd.n22 307.762
R5417 dvdd.n549 dvdd.n15 307.762
R5418 dvdd.t40 dvdd.t42 264.262
R5419 dvdd.t44 dvdd.t40 264.262
R5420 dvdd.t120 dvdd.t44 264.262
R5421 dvdd.t110 dvdd.t120 264.262
R5422 dvdd.t102 dvdd.t110 264.262
R5423 dvdd.t100 dvdd.t102 264.262
R5424 dvdd.t86 dvdd.t100 264.262
R5425 dvdd.t280 dvdd.t86 264.262
R5426 dvdd.t80 dvdd.t280 264.262
R5427 dvdd.t84 dvdd.t80 264.262
R5428 dvdd.t278 dvdd.t84 264.262
R5429 dvdd.t82 dvdd.t278 264.262
R5430 dvdd.n214 dvdd.t25 250.785
R5431 dvdd.n75 dvdd.t144 250.785
R5432 dvdd.n131 dvdd.t321 250.785
R5433 dvdd.n289 dvdd.t267 250.785
R5434 dvdd.n420 dvdd.t219 246.106
R5435 dvdd.n5 dvdd.t7 246.106
R5436 dvdd.n265 dvdd.t105 244.737
R5437 dvdd.n126 dvdd.t176 244.737
R5438 dvdd.n182 dvdd.t69 244.737
R5439 dvdd.n349 dvdd.t53 244.737
R5440 dvdd.n285 dvdd.t229 244.737
R5441 dvdd.n481 dvdd.t122 241.409
R5442 dvdd.n494 dvdd.t117 240.538
R5443 dvdd.n186 dvdd.t119 240.488
R5444 dvdd.n185 dvdd.t83 228.669
R5445 dvdd.t64 dvdd.n502 224.668
R5446 dvdd.t220 dvdd.t58 223.429
R5447 dvdd.t60 dvdd.t220 223.429
R5448 dvdd.t258 dvdd.t248 221.054
R5449 dvdd.t250 dvdd.t258 221.054
R5450 dvdd.t272 dvdd.t250 221.054
R5451 dvdd.t252 dvdd.t272 221.054
R5452 dvdd.t264 dvdd.t252 221.054
R5453 dvdd.t246 dvdd.t264 221.054
R5454 dvdd.t268 dvdd.t246 221.054
R5455 dvdd.t254 dvdd.t268 221.054
R5456 dvdd.t270 dvdd.t254 221.054
R5457 dvdd.t256 dvdd.t270 221.054
R5458 dvdd.t260 dvdd.t256 221.054
R5459 dvdd.t274 dvdd.t260 221.054
R5460 dvdd.t262 dvdd.t276 221.054
R5461 dvdd.t276 dvdd.t266 221.054
R5462 dvdd.t230 dvdd.t226 221.054
R5463 dvdd.t226 dvdd.t232 221.054
R5464 dvdd.t232 dvdd.t228 221.054
R5465 dvdd.t48 dvdd.t50 221.054
R5466 dvdd.t50 dvdd.t46 221.054
R5467 dvdd.t46 dvdd.t52 221.054
R5468 dvdd.t145 dvdd.t165 215.677
R5469 dvdd.t135 dvdd.t145 215.677
R5470 dvdd.t147 dvdd.t135 215.677
R5471 dvdd.t159 dvdd.t147 215.677
R5472 dvdd.t151 dvdd.t159 215.677
R5473 dvdd.t153 dvdd.t151 215.677
R5474 dvdd.t141 dvdd.t153 215.677
R5475 dvdd.t163 dvdd.t141 215.677
R5476 dvdd.t137 dvdd.t163 215.677
R5477 dvdd.t155 dvdd.t137 215.677
R5478 dvdd.t139 dvdd.t157 215.677
R5479 dvdd.t157 dvdd.t149 215.677
R5480 dvdd.t149 dvdd.t161 215.677
R5481 dvdd.t161 dvdd.t143 215.677
R5482 dvdd.t179 dvdd.t177 215.677
R5483 dvdd.t177 dvdd.t181 215.677
R5484 dvdd.t181 dvdd.t175 215.677
R5485 dvdd.t290 dvdd.t310 215.677
R5486 dvdd.t312 dvdd.t290 215.677
R5487 dvdd.t292 dvdd.t312 215.677
R5488 dvdd.t304 dvdd.t292 215.677
R5489 dvdd.t296 dvdd.t304 215.677
R5490 dvdd.t298 dvdd.t296 215.677
R5491 dvdd.t318 dvdd.t298 215.677
R5492 dvdd.t308 dvdd.t318 215.677
R5493 dvdd.t314 dvdd.t308 215.677
R5494 dvdd.t300 dvdd.t314 215.677
R5495 dvdd.t316 dvdd.t302 215.677
R5496 dvdd.t302 dvdd.t294 215.677
R5497 dvdd.t294 dvdd.t306 215.677
R5498 dvdd.t306 dvdd.t320 215.677
R5499 dvdd.t72 dvdd.t66 215.677
R5500 dvdd.t66 dvdd.t70 215.677
R5501 dvdd.t70 dvdd.t68 215.677
R5502 dvdd.t26 dvdd.t14 212.8
R5503 dvdd.t16 dvdd.t26 212.8
R5504 dvdd.t28 dvdd.t16 212.8
R5505 dvdd.t8 dvdd.t28 212.8
R5506 dvdd.t32 dvdd.t8 212.8
R5507 dvdd.t34 dvdd.t32 212.8
R5508 dvdd.t22 dvdd.t34 212.8
R5509 dvdd.t12 dvdd.t22 212.8
R5510 dvdd.t18 dvdd.t12 212.8
R5511 dvdd.t36 dvdd.t18 212.8
R5512 dvdd.t20 dvdd.t38 212.8
R5513 dvdd.t38 dvdd.t30 212.8
R5514 dvdd.t30 dvdd.t10 212.8
R5515 dvdd.t10 dvdd.t24 212.8
R5516 dvdd.t108 dvdd.t106 212.8
R5517 dvdd.t106 dvdd.t112 212.8
R5518 dvdd.t112 dvdd.t104 212.8
R5519 dvdd.n422 dvdd.n415 205.5
R5520 dvdd.n7 dvdd.n0 205.5
R5521 dvdd.t266 dvdd 205.263
R5522 dvdd.n483 dvdd.n477 200.31
R5523 dvdd.n492 dvdd.n489 200.31
R5524 dvdd.n491 dvdd.n490 200.31
R5525 dvdd.n482 dvdd.n478 200.31
R5526 dvdd.n480 dvdd.n479 200.31
R5527 dvdd.n462 dvdd.n461 200.31
R5528 dvdd.t143 dvdd 200.27
R5529 dvdd.t320 dvdd 200.27
R5530 dvdd.n513 dvdd.n512 200.173
R5531 dvdd.n486 dvdd.n485 200.115
R5532 dvdd.n198 dvdd.n197 200.105
R5533 dvdd.n199 dvdd.n196 200.105
R5534 dvdd.n200 dvdd.n195 200.105
R5535 dvdd.n194 dvdd.n189 200.105
R5536 dvdd.n193 dvdd.n190 200.105
R5537 dvdd.n192 dvdd.n191 200.105
R5538 dvdd.n486 dvdd.n484 200.095
R5539 dvdd.n488 dvdd.n487 200.034
R5540 dvdd.t24 dvdd 197.601
R5541 dvdd.t228 dvdd 197.369
R5542 dvdd.t52 dvdd 197.369
R5543 dvdd.t175 dvdd 192.569
R5544 dvdd.t68 dvdd 192.569
R5545 dvdd.t104 dvdd 190
R5546 dvdd.n356 dvdd.n353 185
R5547 dvdd.n357 dvdd.n356 185
R5548 dvdd.n363 dvdd.n360 185
R5549 dvdd.n364 dvdd.n363 185
R5550 dvdd.n370 dvdd.n367 185
R5551 dvdd.n371 dvdd.n370 185
R5552 dvdd.n377 dvdd.n374 185
R5553 dvdd.n378 dvdd.n377 185
R5554 dvdd.n384 dvdd.n381 185
R5555 dvdd.n385 dvdd.n384 185
R5556 dvdd.n391 dvdd.n388 185
R5557 dvdd.n392 dvdd.n391 185
R5558 dvdd.n398 dvdd.n395 185
R5559 dvdd.n399 dvdd.n398 185
R5560 dvdd.n405 dvdd.n402 185
R5561 dvdd.n406 dvdd.n405 185
R5562 dvdd.n412 dvdd.n409 185
R5563 dvdd.n413 dvdd.n412 185
R5564 dvdd.n68 dvdd.n65 185
R5565 dvdd.n69 dvdd.n68 185
R5566 dvdd.n61 dvdd.n58 185
R5567 dvdd.n62 dvdd.n61 185
R5568 dvdd.n54 dvdd.n51 185
R5569 dvdd.n55 dvdd.n54 185
R5570 dvdd.n47 dvdd.n44 185
R5571 dvdd.n48 dvdd.n47 185
R5572 dvdd.n40 dvdd.n37 185
R5573 dvdd.n41 dvdd.n40 185
R5574 dvdd.n33 dvdd.n30 185
R5575 dvdd.n34 dvdd.n33 185
R5576 dvdd.n26 dvdd.n23 185
R5577 dvdd.n27 dvdd.n26 185
R5578 dvdd.n19 dvdd.n16 185
R5579 dvdd.n20 dvdd.n19 185
R5580 dvdd.n12 dvdd.n9 185
R5581 dvdd.n13 dvdd.n12 185
R5582 dvdd.t58 dvdd.t123 180.129
R5583 dvdd.n504 dvdd.t133 175.306
R5584 dvdd.t189 dvdd.n503 174.066
R5585 dvdd.n325 dvdd.t274 171.054
R5586 dvdd.n419 dvdd.t205 157.446
R5587 dvdd.n4 dvdd.t6 157.446
R5588 dvdd.n107 dvdd.t139 146.351
R5589 dvdd.n163 dvdd.t316 146.351
R5590 dvdd.t131 dvdd.t118 145.488
R5591 dvdd.n246 dvdd.t20 141.868
R5592 dvdd.t62 dvdd.t64 136.828
R5593 dvdd.t222 dvdd.t62 136.828
R5594 dvdd.t282 dvdd.t222 136.828
R5595 dvdd.t284 dvdd.t282 136.828
R5596 dvdd.t286 dvdd.t284 136.828
R5597 dvdd.t123 dvdd.t286 136.828
R5598 dvdd.t191 dvdd.t189 136.828
R5599 dvdd.t187 dvdd.t191 136.828
R5600 dvdd.t193 dvdd.t187 136.828
R5601 dvdd.t183 dvdd.t193 136.828
R5602 dvdd.t185 dvdd.t183 136.828
R5603 dvdd.t288 dvdd.n355 129.546
R5604 dvdd.t74 dvdd.n362 129.546
R5605 dvdd.t90 dvdd.n369 129.546
R5606 dvdd.t54 dvdd.n376 129.546
R5607 dvdd.t224 dvdd.n383 129.546
R5608 dvdd.t240 dvdd.n390 129.546
R5609 dvdd.t217 dvdd.n397 129.546
R5610 dvdd.t76 dvdd.n404 129.546
R5611 dvdd.t88 dvdd.n411 129.546
R5612 dvdd.t78 dvdd.n67 129.546
R5613 dvdd.t56 dvdd.n60 129.546
R5614 dvdd.t0 dvdd.n53 129.546
R5615 dvdd.t2 dvdd.n46 129.546
R5616 dvdd.t98 dvdd.n39 129.546
R5617 dvdd.t238 dvdd.n32 129.546
R5618 dvdd.t96 dvdd.n25 129.546
R5619 dvdd.t242 dvdd.n18 129.546
R5620 dvdd.t127 dvdd.n11 129.546
R5621 dvdd.t203 dvdd.n416 127.638
R5622 dvdd.t92 dvdd.n1 127.638
R5623 dvdd.t115 dvdd.t131 117.776
R5624 dvdd.t125 dvdd.t185 109.983
R5625 dvdd.t118 dvdd.t95 109.983
R5626 dvdd.n358 dvdd.n353 101.644
R5627 dvdd.n365 dvdd.n360 101.644
R5628 dvdd.n372 dvdd.n367 101.644
R5629 dvdd.n379 dvdd.n374 101.644
R5630 dvdd.n386 dvdd.n381 101.644
R5631 dvdd.n393 dvdd.n388 101.644
R5632 dvdd.n400 dvdd.n395 101.644
R5633 dvdd.n407 dvdd.n402 101.644
R5634 dvdd.n414 dvdd.n409 101.644
R5635 dvdd.n70 dvdd.n65 101.644
R5636 dvdd.n63 dvdd.n58 101.644
R5637 dvdd.n56 dvdd.n51 101.644
R5638 dvdd.n49 dvdd.n44 101.644
R5639 dvdd.n42 dvdd.n37 101.644
R5640 dvdd.n35 dvdd.n30 101.644
R5641 dvdd.n28 dvdd.n23 101.644
R5642 dvdd.n21 dvdd.n16 101.644
R5643 dvdd.n14 dvdd.n9 101.644
R5644 dvdd.n421 dvdd.n416 95.8438
R5645 dvdd.n6 dvdd.n1 95.8438
R5646 dvdd.n418 dvdd.n417 92.5005
R5647 dvdd.n358 dvdd.n357 92.5005
R5648 dvdd.n365 dvdd.n364 92.5005
R5649 dvdd.n372 dvdd.n371 92.5005
R5650 dvdd.n379 dvdd.n378 92.5005
R5651 dvdd.n386 dvdd.n385 92.5005
R5652 dvdd.n393 dvdd.n392 92.5005
R5653 dvdd.n400 dvdd.n399 92.5005
R5654 dvdd.n407 dvdd.n406 92.5005
R5655 dvdd.n414 dvdd.n413 92.5005
R5656 dvdd.n3 dvdd.n2 92.5005
R5657 dvdd.n70 dvdd.n69 92.5005
R5658 dvdd.n63 dvdd.n62 92.5005
R5659 dvdd.n56 dvdd.n55 92.5005
R5660 dvdd.n49 dvdd.n48 92.5005
R5661 dvdd.n42 dvdd.n41 92.5005
R5662 dvdd.n35 dvdd.n34 92.5005
R5663 dvdd.n28 dvdd.n27 92.5005
R5664 dvdd.n21 dvdd.n20 92.5005
R5665 dvdd.n14 dvdd.n13 92.5005
R5666 dvdd.t95 dvdd.t125 83.1363
R5667 dvdd.n418 dvdd.n416 82.3534
R5668 dvdd.n3 dvdd.n1 82.3534
R5669 dvdd.t133 dvdd.t115 78.8063
R5670 dvdd.n355 dvdd.n354 77.057
R5671 dvdd.n362 dvdd.n361 77.057
R5672 dvdd.n369 dvdd.n368 77.057
R5673 dvdd.n376 dvdd.n375 77.057
R5674 dvdd.n383 dvdd.n382 77.057
R5675 dvdd.n390 dvdd.n389 77.057
R5676 dvdd.n397 dvdd.n396 77.057
R5677 dvdd.n404 dvdd.n403 77.057
R5678 dvdd.n411 dvdd.n410 77.057
R5679 dvdd.n67 dvdd.n66 77.057
R5680 dvdd.n60 dvdd.n59 77.057
R5681 dvdd.n53 dvdd.n52 77.057
R5682 dvdd.n46 dvdd.n45 77.057
R5683 dvdd.n39 dvdd.n38 77.057
R5684 dvdd.n32 dvdd.n31 77.057
R5685 dvdd.n25 dvdd.n24 77.057
R5686 dvdd.n18 dvdd.n17 77.057
R5687 dvdd.n11 dvdd.n10 77.057
R5688 dvdd.n246 dvdd.t36 70.9338
R5689 dvdd.n107 dvdd.t155 69.3248
R5690 dvdd.n163 dvdd.t300 69.3248
R5691 dvdd.n356 dvdd.t288 67.8576
R5692 dvdd.n363 dvdd.t74 67.8576
R5693 dvdd.n370 dvdd.t90 67.8576
R5694 dvdd.n377 dvdd.t54 67.8576
R5695 dvdd.n384 dvdd.t224 67.8576
R5696 dvdd.n391 dvdd.t240 67.8576
R5697 dvdd.n398 dvdd.t217 67.8576
R5698 dvdd.n405 dvdd.t76 67.8576
R5699 dvdd.n412 dvdd.t88 67.8576
R5700 dvdd.n68 dvdd.t78 67.8576
R5701 dvdd.n61 dvdd.t56 67.8576
R5702 dvdd.n54 dvdd.t0 67.8576
R5703 dvdd.n47 dvdd.t2 67.8576
R5704 dvdd.n40 dvdd.t98 67.8576
R5705 dvdd.n33 dvdd.t238 67.8576
R5706 dvdd.n26 dvdd.t96 67.8576
R5707 dvdd.n19 dvdd.t242 67.8576
R5708 dvdd.n12 dvdd.t127 67.8576
R5709 dvdd.n417 dvdd.t203 55.9594
R5710 dvdd.n417 dvdd.t205 55.9594
R5711 dvdd.n2 dvdd.t92 55.9594
R5712 dvdd.n2 dvdd.t6 55.9594
R5713 dvdd.n325 dvdd.t262 50.0005
R5714 dvdd.n355 dvdd.t201 47.2949
R5715 dvdd.n362 dvdd.t199 47.2949
R5716 dvdd.n369 dvdd.t213 47.2949
R5717 dvdd.n376 dvdd.t129 47.2949
R5718 dvdd.n383 dvdd.t236 47.2949
R5719 dvdd.n390 dvdd.t173 47.2949
R5720 dvdd.n397 dvdd.t207 47.2949
R5721 dvdd.n404 dvdd.t171 47.2949
R5722 dvdd.n411 dvdd.t195 47.2949
R5723 dvdd.n67 dvdd.t234 47.2949
R5724 dvdd.n60 dvdd.t211 47.2949
R5725 dvdd.n53 dvdd.t209 47.2949
R5726 dvdd.n46 dvdd.t4 47.2949
R5727 dvdd.n39 dvdd.t244 47.2949
R5728 dvdd.n32 dvdd.t197 47.2949
R5729 dvdd.n25 dvdd.t169 47.2949
R5730 dvdd.n18 dvdd.t215 47.2949
R5731 dvdd.n11 dvdd.t167 47.2949
R5732 dvdd.n206 dvdd.n205 46.2505
R5733 dvdd.n204 dvdd.n187 46.2505
R5734 dvdd.n507 dvdd.n506 45.9299
R5735 dvdd.n420 dvdd.n419 33.4807
R5736 dvdd.n5 dvdd.n4 33.4807
R5737 dvdd.n352 dvdd.t289 32.8338
R5738 dvdd.n352 dvdd.t202 32.8338
R5739 dvdd.n359 dvdd.t75 32.8338
R5740 dvdd.n359 dvdd.t200 32.8338
R5741 dvdd.n366 dvdd.t91 32.8338
R5742 dvdd.n366 dvdd.t214 32.8338
R5743 dvdd.n373 dvdd.t55 32.8338
R5744 dvdd.n373 dvdd.t130 32.8338
R5745 dvdd.n380 dvdd.t225 32.8338
R5746 dvdd.n380 dvdd.t237 32.8338
R5747 dvdd.n387 dvdd.t241 32.8338
R5748 dvdd.n387 dvdd.t174 32.8338
R5749 dvdd.n394 dvdd.t218 32.8338
R5750 dvdd.n394 dvdd.t208 32.8338
R5751 dvdd.n401 dvdd.t77 32.8338
R5752 dvdd.n401 dvdd.t172 32.8338
R5753 dvdd.n408 dvdd.t89 32.8338
R5754 dvdd.n408 dvdd.t196 32.8338
R5755 dvdd.n71 dvdd.t79 32.8338
R5756 dvdd.n71 dvdd.t235 32.8338
R5757 dvdd.n64 dvdd.t57 32.8338
R5758 dvdd.n64 dvdd.t212 32.8338
R5759 dvdd.n57 dvdd.t1 32.8338
R5760 dvdd.n57 dvdd.t210 32.8338
R5761 dvdd.n50 dvdd.t3 32.8338
R5762 dvdd.n50 dvdd.t5 32.8338
R5763 dvdd.n43 dvdd.t99 32.8338
R5764 dvdd.n43 dvdd.t245 32.8338
R5765 dvdd.n36 dvdd.t239 32.8338
R5766 dvdd.n36 dvdd.t198 32.8338
R5767 dvdd.n29 dvdd.t97 32.8338
R5768 dvdd.n29 dvdd.t170 32.8338
R5769 dvdd.n22 dvdd.t243 32.8338
R5770 dvdd.n22 dvdd.t216 32.8338
R5771 dvdd.n15 dvdd.t128 32.8338
R5772 dvdd.n15 dvdd.t168 32.8338
R5773 dvdd.n357 dvdd.n354 30.8889
R5774 dvdd.n354 dvdd.n353 30.8889
R5775 dvdd.n364 dvdd.n361 30.8889
R5776 dvdd.n361 dvdd.n360 30.8889
R5777 dvdd.n371 dvdd.n368 30.8889
R5778 dvdd.n368 dvdd.n367 30.8889
R5779 dvdd.n378 dvdd.n375 30.8889
R5780 dvdd.n375 dvdd.n374 30.8889
R5781 dvdd.n385 dvdd.n382 30.8889
R5782 dvdd.n382 dvdd.n381 30.8889
R5783 dvdd.n392 dvdd.n389 30.8889
R5784 dvdd.n389 dvdd.n388 30.8889
R5785 dvdd.n399 dvdd.n396 30.8889
R5786 dvdd.n396 dvdd.n395 30.8889
R5787 dvdd.n406 dvdd.n403 30.8889
R5788 dvdd.n403 dvdd.n402 30.8889
R5789 dvdd.n413 dvdd.n410 30.8889
R5790 dvdd.n410 dvdd.n409 30.8889
R5791 dvdd.n69 dvdd.n66 30.8889
R5792 dvdd.n66 dvdd.n65 30.8889
R5793 dvdd.n62 dvdd.n59 30.8889
R5794 dvdd.n59 dvdd.n58 30.8889
R5795 dvdd.n55 dvdd.n52 30.8889
R5796 dvdd.n52 dvdd.n51 30.8889
R5797 dvdd.n48 dvdd.n45 30.8889
R5798 dvdd.n45 dvdd.n44 30.8889
R5799 dvdd.n41 dvdd.n38 30.8889
R5800 dvdd.n38 dvdd.n37 30.8889
R5801 dvdd.n34 dvdd.n31 30.8889
R5802 dvdd.n31 dvdd.n30 30.8889
R5803 dvdd.n27 dvdd.n24 30.8889
R5804 dvdd.n24 dvdd.n23 30.8889
R5805 dvdd.n20 dvdd.n17 30.8889
R5806 dvdd.n17 dvdd.n16 30.8889
R5807 dvdd.n13 dvdd.n10 30.8889
R5808 dvdd.n10 dvdd.n9 30.8889
R5809 dvdd.n487 dvdd.t126 29.5505
R5810 dvdd.n514 dvdd.n513 29.3154
R5811 dvdd.n197 dvdd.t85 28.5655
R5812 dvdd.n197 dvdd.t279 28.5655
R5813 dvdd.n196 dvdd.t281 28.5655
R5814 dvdd.n196 dvdd.t81 28.5655
R5815 dvdd.n195 dvdd.t101 28.5655
R5816 dvdd.n195 dvdd.t87 28.5655
R5817 dvdd.n189 dvdd.t111 28.5655
R5818 dvdd.n189 dvdd.t103 28.5655
R5819 dvdd.n190 dvdd.t45 28.5655
R5820 dvdd.n190 dvdd.t121 28.5655
R5821 dvdd.n191 dvdd.t43 28.5655
R5822 dvdd.n191 dvdd.t41 28.5655
R5823 dvdd.n477 dvdd.t61 28.5655
R5824 dvdd.n477 dvdd.t190 28.5655
R5825 dvdd.n485 dvdd.t116 28.5655
R5826 dvdd.n485 dvdd.t134 28.5655
R5827 dvdd.n484 dvdd.t132 28.5655
R5828 dvdd.t116 dvdd.n484 28.5655
R5829 dvdd.n487 dvdd.t186 28.5655
R5830 dvdd.n489 dvdd.t194 28.5655
R5831 dvdd.n489 dvdd.t184 28.5655
R5832 dvdd.n490 dvdd.t192 28.5655
R5833 dvdd.n490 dvdd.t188 28.5655
R5834 dvdd.n478 dvdd.t59 28.5655
R5835 dvdd.n478 dvdd.t221 28.5655
R5836 dvdd.n479 dvdd.t285 28.5655
R5837 dvdd.n479 dvdd.t287 28.5655
R5838 dvdd.n461 dvdd.t223 28.5655
R5839 dvdd.n461 dvdd.t283 28.5655
R5840 dvdd.n512 dvdd.t65 28.5655
R5841 dvdd.n512 dvdd.t63 28.5655
R5842 dvdd.n419 dvdd.n418 27.7986
R5843 dvdd.n4 dvdd.n3 27.7986
R5844 dvdd.n212 dvdd.t107 26.5955
R5845 dvdd.n212 dvdd.t113 26.5955
R5846 dvdd.n216 dvdd.t31 26.5955
R5847 dvdd.n216 dvdd.t11 26.5955
R5848 dvdd.n217 dvdd.t21 26.5955
R5849 dvdd.n217 dvdd.t39 26.5955
R5850 dvdd.n220 dvdd.t19 26.5955
R5851 dvdd.n220 dvdd.t37 26.5955
R5852 dvdd.n237 dvdd.t23 26.5955
R5853 dvdd.n237 dvdd.t13 26.5955
R5854 dvdd.n223 dvdd.t33 26.5955
R5855 dvdd.n223 dvdd.t35 26.5955
R5856 dvdd.n228 dvdd.t29 26.5955
R5857 dvdd.n228 dvdd.t9 26.5955
R5858 dvdd.n226 dvdd.t27 26.5955
R5859 dvdd.n226 dvdd.t17 26.5955
R5860 dvdd.n73 dvdd.t178 26.5955
R5861 dvdd.n73 dvdd.t182 26.5955
R5862 dvdd.n77 dvdd.t150 26.5955
R5863 dvdd.n77 dvdd.t162 26.5955
R5864 dvdd.n78 dvdd.t140 26.5955
R5865 dvdd.n78 dvdd.t158 26.5955
R5866 dvdd.n81 dvdd.t138 26.5955
R5867 dvdd.n81 dvdd.t156 26.5955
R5868 dvdd.n98 dvdd.t142 26.5955
R5869 dvdd.n98 dvdd.t164 26.5955
R5870 dvdd.n84 dvdd.t152 26.5955
R5871 dvdd.n84 dvdd.t154 26.5955
R5872 dvdd.n89 dvdd.t148 26.5955
R5873 dvdd.n89 dvdd.t160 26.5955
R5874 dvdd.n87 dvdd.t146 26.5955
R5875 dvdd.n87 dvdd.t136 26.5955
R5876 dvdd.n129 dvdd.t67 26.5955
R5877 dvdd.n129 dvdd.t71 26.5955
R5878 dvdd.n133 dvdd.t295 26.5955
R5879 dvdd.n133 dvdd.t307 26.5955
R5880 dvdd.n134 dvdd.t317 26.5955
R5881 dvdd.n134 dvdd.t303 26.5955
R5882 dvdd.n137 dvdd.t315 26.5955
R5883 dvdd.n137 dvdd.t301 26.5955
R5884 dvdd.n154 dvdd.t319 26.5955
R5885 dvdd.n154 dvdd.t309 26.5955
R5886 dvdd.n140 dvdd.t297 26.5955
R5887 dvdd.n140 dvdd.t299 26.5955
R5888 dvdd.n145 dvdd.t293 26.5955
R5889 dvdd.n145 dvdd.t305 26.5955
R5890 dvdd.n143 dvdd.t291 26.5955
R5891 dvdd.n143 dvdd.t313 26.5955
R5892 dvdd.n287 dvdd.t227 26.5955
R5893 dvdd.n287 dvdd.t233 26.5955
R5894 dvdd.n283 dvdd.t51 26.5955
R5895 dvdd.n283 dvdd.t47 26.5955
R5896 dvdd.n291 dvdd.t263 26.5955
R5897 dvdd.n291 dvdd.t277 26.5955
R5898 dvdd.n292 dvdd.t261 26.5955
R5899 dvdd.n292 dvdd.t275 26.5955
R5900 dvdd.n295 dvdd.t271 26.5955
R5901 dvdd.n295 dvdd.t257 26.5955
R5902 dvdd.n312 dvdd.t269 26.5955
R5903 dvdd.n312 dvdd.t255 26.5955
R5904 dvdd.n298 dvdd.t265 26.5955
R5905 dvdd.n298 dvdd.t247 26.5955
R5906 dvdd.n303 dvdd.t273 26.5955
R5907 dvdd.n303 dvdd.t253 26.5955
R5908 dvdd.n301 dvdd.t259 26.5955
R5909 dvdd.n301 dvdd.t251 26.5955
R5910 dvdd.n415 dvdd.t204 24.6255
R5911 dvdd.n415 dvdd.t206 24.6255
R5912 dvdd.n0 dvdd.t93 24.6255
R5913 dvdd.n0 dvdd.t94 24.6255
R5914 dvdd.n457 dvdd.n456 22.5272
R5915 dvdd.n453 dvdd.n452 22.5272
R5916 dvdd.n449 dvdd.n448 22.5272
R5917 dvdd.n445 dvdd.n444 22.5272
R5918 dvdd.n441 dvdd.n440 22.5272
R5919 dvdd.n437 dvdd.n436 22.5272
R5920 dvdd.n433 dvdd.n432 22.5272
R5921 dvdd.n429 dvdd.n428 22.5272
R5922 dvdd.n425 dvdd.n424 22.5272
R5923 dvdd.n519 dvdd.n518 22.5272
R5924 dvdd.n523 dvdd.n522 22.5272
R5925 dvdd.n527 dvdd.n526 22.5272
R5926 dvdd.n531 dvdd.n530 22.5272
R5927 dvdd.n535 dvdd.n534 22.5272
R5928 dvdd.n539 dvdd.n538 22.5272
R5929 dvdd.n543 dvdd.n542 22.5272
R5930 dvdd.n547 dvdd.n546 22.5272
R5931 dvdd.n551 dvdd.n550 22.5272
R5932 dvdd.n476 dvdd.n475 18.9204
R5933 dvdd.n309 dvdd.n299 18.1174
R5934 dvdd.n314 dvdd.n311 18.1174
R5935 dvdd.n318 dvdd.n296 18.1174
R5936 dvdd.n321 dvdd.n320 18.1174
R5937 dvdd.n329 dvdd.n328 18.1174
R5938 dvdd.n333 dvdd.n332 18.1174
R5939 dvdd.n337 dvdd.n336 18.1174
R5940 dvdd.n338 dvdd.n337 18.1174
R5941 dvdd.n343 dvdd.n341 18.1174
R5942 dvdd.n347 dvdd.n284 18.1174
R5943 dvdd.n348 dvdd.n347 18.1174
R5944 dvdd.n305 dvdd.n302 17.9205
R5945 dvdd.n458 dvdd.n457 17.4938
R5946 dvdd.n454 dvdd.n453 17.4938
R5947 dvdd.n450 dvdd.n449 17.4938
R5948 dvdd.n446 dvdd.n445 17.4938
R5949 dvdd.n442 dvdd.n441 17.4938
R5950 dvdd.n438 dvdd.n437 17.4938
R5951 dvdd.n434 dvdd.n433 17.4938
R5952 dvdd.n430 dvdd.n429 17.4938
R5953 dvdd.n426 dvdd.n425 17.4938
R5954 dvdd.n518 dvdd.n517 17.4938
R5955 dvdd.n522 dvdd.n521 17.4938
R5956 dvdd.n526 dvdd.n525 17.4938
R5957 dvdd.n530 dvdd.n529 17.4938
R5958 dvdd.n534 dvdd.n533 17.4938
R5959 dvdd.n538 dvdd.n537 17.4938
R5960 dvdd.n542 dvdd.n541 17.4938
R5961 dvdd.n546 dvdd.n545 17.4938
R5962 dvdd.n550 dvdd.n549 17.4938
R5963 dvdd.n338 dvdd.n285 16.9359
R5964 dvdd.n349 dvdd.n348 16.9359
R5965 dvdd.n234 dvdd.n224 16.132
R5966 dvdd.n239 dvdd.n236 16.132
R5967 dvdd.n243 dvdd.n221 16.132
R5968 dvdd.n254 dvdd.n253 16.132
R5969 dvdd.n259 dvdd.n257 16.132
R5970 dvdd.n263 dvdd.n213 16.132
R5971 dvdd.n264 dvdd.n263 16.132
R5972 dvdd.n230 dvdd.n227 15.9567
R5973 dvdd.n95 dvdd.n85 15.914
R5974 dvdd.n100 dvdd.n97 15.914
R5975 dvdd.n104 dvdd.n82 15.914
R5976 dvdd.n115 dvdd.n114 15.914
R5977 dvdd.n120 dvdd.n118 15.914
R5978 dvdd.n124 dvdd.n74 15.914
R5979 dvdd.n125 dvdd.n124 15.914
R5980 dvdd.n151 dvdd.n141 15.914
R5981 dvdd.n156 dvdd.n153 15.914
R5982 dvdd.n160 dvdd.n138 15.914
R5983 dvdd.n171 dvdd.n170 15.914
R5984 dvdd.n176 dvdd.n174 15.914
R5985 dvdd.n180 dvdd.n130 15.914
R5986 dvdd.n181 dvdd.n180 15.914
R5987 dvdd.n336 dvdd.n288 15.7543
R5988 dvdd.n342 dvdd.n284 15.7543
R5989 dvdd.n91 dvdd.n88 15.741
R5990 dvdd.n147 dvdd.n144 15.741
R5991 dvdd.n252 dvdd.n251 15.606
R5992 dvdd.n324 dvdd.n293 15.5574
R5993 dvdd.n421 dvdd 15.5495
R5994 dvdd.n6 dvdd 15.5495
R5995 dvdd.n113 dvdd.n112 15.3951
R5996 dvdd.n169 dvdd.n168 15.3951
R5997 dvdd.n305 dvdd.n304 15.1636
R5998 dvdd.n329 dvdd.n289 15.1636
R5999 dvdd.n265 dvdd.n264 15.08
R6000 dvdd.n248 dvdd.n247 14.9046
R6001 dvdd.n109 dvdd.n108 14.8762
R6002 dvdd.n126 dvdd.n125 14.8762
R6003 dvdd.n165 dvdd.n164 14.8762
R6004 dvdd.n182 dvdd.n181 14.8762
R6005 dvdd.n247 dvdd.n246 14.2313
R6006 dvdd.n505 dvdd.n504 14.2313
R6007 dvdd.n502 dvdd.n498 14.2313
R6008 dvdd.n258 dvdd.n213 14.0279
R6009 dvdd.n251 dvdd.n218 13.8526
R6010 dvdd.n119 dvdd.n74 13.8383
R6011 dvdd.n175 dvdd.n130 13.8383
R6012 dvdd.n108 dvdd.n107 13.7042
R6013 dvdd.n164 dvdd.n163 13.7042
R6014 dvdd.n112 dvdd.n79 13.6654
R6015 dvdd.n168 dvdd.n135 13.6654
R6016 dvdd.n230 dvdd.n229 13.5019
R6017 dvdd.n254 dvdd.n214 13.5019
R6018 dvdd.n91 dvdd.n90 13.3194
R6019 dvdd.n115 dvdd.n75 13.3194
R6020 dvdd.n147 dvdd.n146 13.3194
R6021 dvdd.n171 dvdd.n131 13.3194
R6022 dvdd.n320 dvdd.n319 12.4067
R6023 dvdd.n310 dvdd.n309 12.0128
R6024 dvdd.n327 dvdd.n326 12.0128
R6025 dvdd.n326 dvdd.n325 11.2126
R6026 dvdd.n245 dvdd.n244 11.0471
R6027 dvdd.n106 dvdd.n105 10.8978
R6028 dvdd.n162 dvdd.n161 10.8978
R6029 dvdd.n235 dvdd.n234 10.6964
R6030 dvdd.n96 dvdd.n95 10.5519
R6031 dvdd.n152 dvdd.n151 10.5519
R6032 dvdd.n350 dvdd.n349 10.482
R6033 dvdd.n266 dvdd.n265 10.3526
R6034 dvdd.n127 dvdd.n126 10.3383
R6035 dvdd.n183 dvdd.n182 10.3383
R6036 dvdd.n423 dvdd.n422 10.0534
R6037 dvdd.n8 dvdd.n7 10.0534
R6038 dvdd.n460 dvdd.n351 9.76224
R6039 dvdd.n279 dvdd.n278 9.50994
R6040 dvdd.n231 dvdd.n230 9.3005
R6041 dvdd.n232 dvdd.n224 9.3005
R6042 dvdd.n234 dvdd.n233 9.3005
R6043 dvdd.n236 dvdd.n222 9.3005
R6044 dvdd.n240 dvdd.n239 9.3005
R6045 dvdd.n241 dvdd.n221 9.3005
R6046 dvdd.n243 dvdd.n242 9.3005
R6047 dvdd.n245 dvdd.n219 9.3005
R6048 dvdd.n249 dvdd.n248 9.3005
R6049 dvdd.n251 dvdd.n250 9.3005
R6050 dvdd.n253 dvdd.n215 9.3005
R6051 dvdd.n255 dvdd.n254 9.3005
R6052 dvdd.n257 dvdd.n256 9.3005
R6053 dvdd.n260 dvdd.n259 9.3005
R6054 dvdd.n261 dvdd.n213 9.3005
R6055 dvdd.n263 dvdd.n262 9.3005
R6056 dvdd.n264 dvdd.n211 9.3005
R6057 dvdd.n125 dvdd.n72 9.3005
R6058 dvdd.n124 dvdd.n123 9.3005
R6059 dvdd.n122 dvdd.n74 9.3005
R6060 dvdd.n121 dvdd.n120 9.3005
R6061 dvdd.n118 dvdd.n117 9.3005
R6062 dvdd.n116 dvdd.n115 9.3005
R6063 dvdd.n114 dvdd.n76 9.3005
R6064 dvdd.n112 dvdd.n111 9.3005
R6065 dvdd.n110 dvdd.n109 9.3005
R6066 dvdd.n106 dvdd.n80 9.3005
R6067 dvdd.n104 dvdd.n103 9.3005
R6068 dvdd.n102 dvdd.n82 9.3005
R6069 dvdd.n101 dvdd.n100 9.3005
R6070 dvdd.n97 dvdd.n83 9.3005
R6071 dvdd.n95 dvdd.n94 9.3005
R6072 dvdd.n93 dvdd.n85 9.3005
R6073 dvdd.n92 dvdd.n91 9.3005
R6074 dvdd.n181 dvdd.n128 9.3005
R6075 dvdd.n180 dvdd.n179 9.3005
R6076 dvdd.n178 dvdd.n130 9.3005
R6077 dvdd.n177 dvdd.n176 9.3005
R6078 dvdd.n174 dvdd.n173 9.3005
R6079 dvdd.n172 dvdd.n171 9.3005
R6080 dvdd.n170 dvdd.n132 9.3005
R6081 dvdd.n168 dvdd.n167 9.3005
R6082 dvdd.n166 dvdd.n165 9.3005
R6083 dvdd.n162 dvdd.n136 9.3005
R6084 dvdd.n160 dvdd.n159 9.3005
R6085 dvdd.n158 dvdd.n138 9.3005
R6086 dvdd.n157 dvdd.n156 9.3005
R6087 dvdd.n153 dvdd.n139 9.3005
R6088 dvdd.n151 dvdd.n150 9.3005
R6089 dvdd.n149 dvdd.n141 9.3005
R6090 dvdd.n148 dvdd.n147 9.3005
R6091 dvdd.n341 dvdd.n340 9.3005
R6092 dvdd.n348 dvdd.n282 9.3005
R6093 dvdd.n347 dvdd.n346 9.3005
R6094 dvdd.n345 dvdd.n284 9.3005
R6095 dvdd.n344 dvdd.n343 9.3005
R6096 dvdd.n339 dvdd.n338 9.3005
R6097 dvdd.n337 dvdd.n286 9.3005
R6098 dvdd.n336 dvdd.n335 9.3005
R6099 dvdd.n334 dvdd.n333 9.3005
R6100 dvdd.n332 dvdd.n331 9.3005
R6101 dvdd.n330 dvdd.n329 9.3005
R6102 dvdd.n328 dvdd.n290 9.3005
R6103 dvdd.n324 dvdd.n323 9.3005
R6104 dvdd.n322 dvdd.n321 9.3005
R6105 dvdd.n320 dvdd.n294 9.3005
R6106 dvdd.n318 dvdd.n317 9.3005
R6107 dvdd.n316 dvdd.n296 9.3005
R6108 dvdd.n315 dvdd.n314 9.3005
R6109 dvdd.n311 dvdd.n297 9.3005
R6110 dvdd.n309 dvdd.n308 9.3005
R6111 dvdd.n307 dvdd.n299 9.3005
R6112 dvdd.n306 dvdd.n305 9.3005
R6113 dvdd.n427 dvdd.n426 9.3005
R6114 dvdd.n431 dvdd.n430 9.3005
R6115 dvdd.n435 dvdd.n434 9.3005
R6116 dvdd.n439 dvdd.n438 9.3005
R6117 dvdd.n443 dvdd.n442 9.3005
R6118 dvdd.n447 dvdd.n446 9.3005
R6119 dvdd.n451 dvdd.n450 9.3005
R6120 dvdd.n455 dvdd.n454 9.3005
R6121 dvdd.n459 dvdd.n458 9.3005
R6122 dvdd.n549 dvdd.n548 9.3005
R6123 dvdd.n545 dvdd.n544 9.3005
R6124 dvdd.n541 dvdd.n540 9.3005
R6125 dvdd.n537 dvdd.n536 9.3005
R6126 dvdd.n533 dvdd.n532 9.3005
R6127 dvdd.n529 dvdd.n528 9.3005
R6128 dvdd.n525 dvdd.n524 9.3005
R6129 dvdd.n521 dvdd.n520 9.3005
R6130 dvdd.n517 dvdd.n516 9.3005
R6131 dvdd.n506 dvdd.n497 9.3005
R6132 dvdd.n313 dvdd.n296 9.25588
R6133 dvdd.n314 dvdd.n313 8.86204
R6134 dvdd.n238 dvdd.n221 8.2416
R6135 dvdd.n99 dvdd.n82 8.13023
R6136 dvdd.n155 dvdd.n138 8.13023
R6137 dvdd.n239 dvdd.n238 7.89091
R6138 dvdd.n100 dvdd.n99 7.78428
R6139 dvdd.n156 dvdd.n155 7.78428
R6140 dvdd.n476 dvdd.n464 7.68556
R6141 dvdd.n422 dvdd.n421 6.58874
R6142 dvdd.n7 dvdd.n6 6.58874
R6143 dvdd.n509 dvdd.n476 6.50028
R6144 dvdd.n302 dvdd.n300 6.14225
R6145 dvdd.n311 dvdd.n310 6.10512
R6146 dvdd.n503 dvdd.t60 6.06249
R6147 dvdd.n207 dvdd.n188 5.96824
R6148 dvdd.t100 dvdd.n188 5.96824
R6149 dvdd.n203 dvdd.n202 5.96824
R6150 dvdd.t100 dvdd.n203 5.96824
R6151 dvdd.n184 dvdd 5.94484
R6152 dvdd.n510 dvdd.n463 5.9447
R6153 dvdd.n496 dvdd.n463 5.94023
R6154 dvdd.n227 dvdd.n225 5.87299
R6155 dvdd.n88 dvdd.n86 5.84114
R6156 dvdd.n144 dvdd.n142 5.84114
R6157 dvdd.n319 dvdd.n318 5.71127
R6158 dvdd.n326 dvdd.n324 5.51435
R6159 dvdd.n236 dvdd.n235 5.43612
R6160 dvdd.n97 dvdd.n96 5.36266
R6161 dvdd.n153 dvdd.n152 5.36266
R6162 dvdd.n351 dvdd 5.14764
R6163 dvdd.n184 dvdd 5.14243
R6164 dvdd.n244 dvdd.n243 5.08543
R6165 dvdd.n105 dvdd.n104 5.01672
R6166 dvdd.n161 dvdd.n160 5.01672
R6167 dvdd.n281 dvdd.n280 4.5005
R6168 dvdd.n457 dvdd.n358 4.32258
R6169 dvdd.n453 dvdd.n365 4.32258
R6170 dvdd.n449 dvdd.n372 4.32258
R6171 dvdd.n445 dvdd.n379 4.32258
R6172 dvdd.n441 dvdd.n386 4.32258
R6173 dvdd.n437 dvdd.n393 4.32258
R6174 dvdd.n433 dvdd.n400 4.32258
R6175 dvdd.n429 dvdd.n407 4.32258
R6176 dvdd.n425 dvdd.n414 4.32258
R6177 dvdd.n518 dvdd.n70 4.32258
R6178 dvdd.n522 dvdd.n63 4.32258
R6179 dvdd.n526 dvdd.n56 4.32258
R6180 dvdd.n530 dvdd.n49 4.32258
R6181 dvdd.n534 dvdd.n42 4.32258
R6182 dvdd.n538 dvdd.n35 4.32258
R6183 dvdd.n542 dvdd.n28 4.32258
R6184 dvdd.n546 dvdd.n21 4.32258
R6185 dvdd.n550 dvdd.n14 4.32258
R6186 dvdd.n509 dvdd.n508 4.29291
R6187 dvdd.n497 dvdd.n496 4.26836
R6188 dvdd.n514 dvdd 4.0955
R6189 dvdd.n460 dvdd 3.73954
R6190 dvdd dvdd.n515 3.73954
R6191 dvdd.n501 dvdd.n500 3.36414
R6192 dvdd.n503 dvdd.n501 3.36414
R6193 dvdd.n507 dvdd.n499 3.36414
R6194 dvdd.n503 dvdd.n499 3.36414
R6195 dvdd.n209 dvdd.n208 3.36211
R6196 dvdd.n421 dvdd.n420 3.34378
R6197 dvdd.n6 dvdd.n5 3.34378
R6198 dvdd.n272 dvdd.n268 3.13609
R6199 dvdd.n273 dvdd.n272 3.13609
R6200 dvdd.n277 dvdd.n276 3.13609
R6201 dvdd.n276 dvdd.n275 3.13609
R6202 dvdd.n304 dvdd.n299 2.95435
R6203 dvdd.n332 dvdd.n289 2.95435
R6204 dvdd.n424 dvdd 2.9391
R6205 dvdd.n428 dvdd 2.9391
R6206 dvdd.n432 dvdd 2.9391
R6207 dvdd.n436 dvdd 2.9391
R6208 dvdd.n440 dvdd 2.9391
R6209 dvdd.n444 dvdd 2.9391
R6210 dvdd.n448 dvdd 2.9391
R6211 dvdd.n452 dvdd 2.9391
R6212 dvdd.n456 dvdd 2.9391
R6213 dvdd dvdd.n547 2.9391
R6214 dvdd dvdd.n543 2.9391
R6215 dvdd dvdd.n539 2.9391
R6216 dvdd dvdd.n535 2.9391
R6217 dvdd dvdd.n531 2.9391
R6218 dvdd dvdd.n527 2.9391
R6219 dvdd dvdd.n523 2.9391
R6220 dvdd dvdd.n519 2.9391
R6221 dvdd dvdd.n551 2.9369
R6222 dvdd.n192 dvdd.n186 2.90005
R6223 dvdd.n469 dvdd.n465 2.80353
R6224 dvdd.n470 dvdd.n469 2.80353
R6225 dvdd.n474 dvdd.n473 2.80353
R6226 dvdd.n473 dvdd.n472 2.80353
R6227 dvdd.n229 dvdd.n224 2.63064
R6228 dvdd.n257 dvdd.n214 2.63064
R6229 dvdd.n90 dvdd.n85 2.59509
R6230 dvdd.n118 dvdd.n75 2.59509
R6231 dvdd.n146 dvdd.n141 2.59509
R6232 dvdd.n174 dvdd.n131 2.59509
R6233 dvdd.n321 dvdd.n293 2.5605
R6234 dvdd.n210 dvdd.n209 2.52884
R6235 dvdd.n333 dvdd.n288 2.36358
R6236 dvdd.n343 dvdd.n342 2.36358
R6237 dvdd.n248 dvdd.n218 2.27995
R6238 dvdd.n109 dvdd.n79 2.24915
R6239 dvdd.n165 dvdd.n135 2.24915
R6240 dvdd.n259 dvdd.n258 2.10461
R6241 dvdd.n120 dvdd.n119 2.07618
R6242 dvdd.n176 dvdd.n175 2.07618
R6243 dvdd.n279 dvdd.n267 1.83443
R6244 dvdd.n280 dvdd.n279 1.72468
R6245 dvdd.n515 dvdd.n460 1.69386
R6246 dvdd.n270 dvdd.n267 1.37087
R6247 dvdd.n274 dvdd.n270 1.37087
R6248 dvdd.n278 dvdd.n269 1.37087
R6249 dvdd.n271 dvdd.n269 1.37087
R6250 dvdd.n281 dvdd.n210 1.26417
R6251 dvdd.n247 dvdd.n245 1.2279
R6252 dvdd.n341 dvdd.n285 1.18204
R6253 dvdd.n92 dvdd.n86 1.06234
R6254 dvdd.n148 dvdd.n142 1.06234
R6255 dvdd.n231 dvdd.n225 1.05227
R6256 dvdd.n108 dvdd.n106 1.03834
R6257 dvdd.n164 dvdd.n162 1.03834
R6258 dvdd.n306 dvdd.n300 0.968765
R6259 dvdd.n208 dvdd.n186 0.955857
R6260 dvdd.n515 dvdd.n514 0.951672
R6261 dvdd.n210 dvdd.n184 0.836438
R6262 dvdd.n483 dvdd.n482 0.787085
R6263 dvdd.n193 dvdd.n192 0.705857
R6264 dvdd.n194 dvdd.n193 0.705857
R6265 dvdd.n200 dvdd.n199 0.705857
R6266 dvdd.n199 dvdd.n198 0.705857
R6267 dvdd.n198 dvdd.n185 0.705857
R6268 dvdd.n351 dvdd.n281 0.691906
R6269 dvdd.n280 dvdd 0.645031
R6270 dvdd.n328 dvdd.n327 0.591269
R6271 dvdd.n201 dvdd.n194 0.529518
R6272 dvdd.n253 dvdd.n252 0.526527
R6273 dvdd.n114 dvdd.n113 0.519419
R6274 dvdd.n170 dvdd.n169 0.519419
R6275 dvdd.n482 dvdd.n481 0.514219
R6276 dvdd.n495 dvdd.n494 0.492878
R6277 dvdd.n480 dvdd.n462 0.482207
R6278 dvdd.n491 dvdd.n483 0.482207
R6279 dvdd.n492 dvdd.n491 0.482207
R6280 dvdd.n493 dvdd.n492 0.482207
R6281 dvdd.n467 dvdd.n464 0.468854
R6282 dvdd.n468 dvdd.n467 0.468854
R6283 dvdd.n475 dvdd.n466 0.468854
R6284 dvdd.n471 dvdd.n466 0.468854
R6285 dvdd.n511 dvdd.n462 0.447146
R6286 dvdd.n496 dvdd.n495 0.419707
R6287 dvdd.n494 dvdd.n493 0.386171
R6288 dvdd.n511 dvdd.n510 0.372451
R6289 dvdd.n481 dvdd.n480 0.361781
R6290 dvdd.n209 dvdd.n185 0.346482
R6291 dvdd.n202 dvdd.n201 0.3105
R6292 dvdd.n208 dvdd.n207 0.3105
R6293 dvdd.n497 dvdd.n483 0.307565
R6294 dvdd.n508 dvdd.n497 0.272821
R6295 dvdd.n510 dvdd.n509 0.252732
R6296 dvdd.n495 dvdd.n486 0.206229
R6297 dvdd.n500 dvdd.n463 0.179346
R6298 dvdd.n508 dvdd.n507 0.179346
R6299 dvdd.n201 dvdd.n200 0.176839
R6300 dvdd.n493 dvdd.n488 0.152674
R6301 dvdd.n423 dvdd 0.121114
R6302 dvdd.n427 dvdd 0.121114
R6303 dvdd.n431 dvdd 0.121114
R6304 dvdd.n435 dvdd 0.121114
R6305 dvdd.n439 dvdd 0.121114
R6306 dvdd.n443 dvdd 0.121114
R6307 dvdd.n447 dvdd 0.121114
R6308 dvdd.n451 dvdd 0.121114
R6309 dvdd.n455 dvdd 0.121114
R6310 dvdd.n459 dvdd 0.121114
R6311 dvdd.n8 dvdd 0.121114
R6312 dvdd.n548 dvdd 0.121114
R6313 dvdd.n544 dvdd 0.121114
R6314 dvdd.n540 dvdd 0.121114
R6315 dvdd.n536 dvdd 0.121114
R6316 dvdd.n532 dvdd 0.121114
R6317 dvdd.n528 dvdd 0.121114
R6318 dvdd.n524 dvdd 0.121114
R6319 dvdd.n520 dvdd 0.121114
R6320 dvdd.n516 dvdd 0.121114
R6321 dvdd.n232 dvdd.n231 0.120292
R6322 dvdd.n233 dvdd.n232 0.120292
R6323 dvdd.n233 dvdd.n222 0.120292
R6324 dvdd.n240 dvdd.n222 0.120292
R6325 dvdd.n241 dvdd.n240 0.120292
R6326 dvdd.n242 dvdd.n241 0.120292
R6327 dvdd.n242 dvdd.n219 0.120292
R6328 dvdd.n249 dvdd.n219 0.120292
R6329 dvdd.n250 dvdd.n249 0.120292
R6330 dvdd.n250 dvdd.n215 0.120292
R6331 dvdd.n255 dvdd.n215 0.120292
R6332 dvdd.n256 dvdd.n255 0.120292
R6333 dvdd.n261 dvdd.n260 0.120292
R6334 dvdd.n262 dvdd.n261 0.120292
R6335 dvdd.n262 dvdd.n211 0.120292
R6336 dvdd.n266 dvdd.n211 0.120292
R6337 dvdd.n93 dvdd.n92 0.120292
R6338 dvdd.n94 dvdd.n93 0.120292
R6339 dvdd.n94 dvdd.n83 0.120292
R6340 dvdd.n101 dvdd.n83 0.120292
R6341 dvdd.n102 dvdd.n101 0.120292
R6342 dvdd.n103 dvdd.n102 0.120292
R6343 dvdd.n103 dvdd.n80 0.120292
R6344 dvdd.n110 dvdd.n80 0.120292
R6345 dvdd.n111 dvdd.n110 0.120292
R6346 dvdd.n111 dvdd.n76 0.120292
R6347 dvdd.n116 dvdd.n76 0.120292
R6348 dvdd.n117 dvdd.n116 0.120292
R6349 dvdd.n122 dvdd.n121 0.120292
R6350 dvdd.n123 dvdd.n122 0.120292
R6351 dvdd.n123 dvdd.n72 0.120292
R6352 dvdd.n127 dvdd.n72 0.120292
R6353 dvdd.n149 dvdd.n148 0.120292
R6354 dvdd.n150 dvdd.n149 0.120292
R6355 dvdd.n150 dvdd.n139 0.120292
R6356 dvdd.n157 dvdd.n139 0.120292
R6357 dvdd.n158 dvdd.n157 0.120292
R6358 dvdd.n159 dvdd.n158 0.120292
R6359 dvdd.n159 dvdd.n136 0.120292
R6360 dvdd.n166 dvdd.n136 0.120292
R6361 dvdd.n167 dvdd.n166 0.120292
R6362 dvdd.n167 dvdd.n132 0.120292
R6363 dvdd.n172 dvdd.n132 0.120292
R6364 dvdd.n173 dvdd.n172 0.120292
R6365 dvdd.n178 dvdd.n177 0.120292
R6366 dvdd.n179 dvdd.n178 0.120292
R6367 dvdd.n179 dvdd.n128 0.120292
R6368 dvdd.n183 dvdd.n128 0.120292
R6369 dvdd.n307 dvdd.n306 0.120292
R6370 dvdd.n308 dvdd.n307 0.120292
R6371 dvdd.n308 dvdd.n297 0.120292
R6372 dvdd.n315 dvdd.n297 0.120292
R6373 dvdd.n316 dvdd.n315 0.120292
R6374 dvdd.n317 dvdd.n316 0.120292
R6375 dvdd.n317 dvdd.n294 0.120292
R6376 dvdd.n322 dvdd.n294 0.120292
R6377 dvdd.n323 dvdd.n322 0.120292
R6378 dvdd.n323 dvdd.n290 0.120292
R6379 dvdd.n330 dvdd.n290 0.120292
R6380 dvdd.n331 dvdd.n330 0.120292
R6381 dvdd.n335 dvdd.n334 0.120292
R6382 dvdd.n335 dvdd.n286 0.120292
R6383 dvdd.n339 dvdd.n286 0.120292
R6384 dvdd.n340 dvdd.n339 0.120292
R6385 dvdd.n345 dvdd.n344 0.120292
R6386 dvdd.n346 dvdd.n345 0.120292
R6387 dvdd.n346 dvdd.n282 0.120292
R6388 dvdd.n350 dvdd.n282 0.120292
R6389 dvdd.n513 dvdd.n511 0.0789314
R6390 dvdd.n260 dvdd 0.0603958
R6391 dvdd.n121 dvdd 0.0603958
R6392 dvdd.n177 dvdd 0.0603958
R6393 dvdd.n334 dvdd 0.0603958
R6394 dvdd.n344 dvdd 0.0603958
R6395 dvdd dvdd.n423 0.0377807
R6396 dvdd.n424 dvdd 0.0377807
R6397 dvdd dvdd.n427 0.0377807
R6398 dvdd.n428 dvdd 0.0377807
R6399 dvdd dvdd.n431 0.0377807
R6400 dvdd.n432 dvdd 0.0377807
R6401 dvdd dvdd.n435 0.0377807
R6402 dvdd.n436 dvdd 0.0377807
R6403 dvdd dvdd.n439 0.0377807
R6404 dvdd.n440 dvdd 0.0377807
R6405 dvdd dvdd.n443 0.0377807
R6406 dvdd.n444 dvdd 0.0377807
R6407 dvdd dvdd.n447 0.0377807
R6408 dvdd.n448 dvdd 0.0377807
R6409 dvdd dvdd.n451 0.0377807
R6410 dvdd.n452 dvdd 0.0377807
R6411 dvdd dvdd.n455 0.0377807
R6412 dvdd.n456 dvdd 0.0377807
R6413 dvdd dvdd.n459 0.0377807
R6414 dvdd dvdd.n8 0.0377807
R6415 dvdd.n551 dvdd 0.0377807
R6416 dvdd.n548 dvdd 0.0377807
R6417 dvdd.n547 dvdd 0.0377807
R6418 dvdd.n544 dvdd 0.0377807
R6419 dvdd.n543 dvdd 0.0377807
R6420 dvdd.n540 dvdd 0.0377807
R6421 dvdd.n539 dvdd 0.0377807
R6422 dvdd.n536 dvdd 0.0377807
R6423 dvdd.n535 dvdd 0.0377807
R6424 dvdd.n532 dvdd 0.0377807
R6425 dvdd.n531 dvdd 0.0377807
R6426 dvdd.n528 dvdd 0.0377807
R6427 dvdd.n527 dvdd 0.0377807
R6428 dvdd.n524 dvdd 0.0377807
R6429 dvdd.n523 dvdd 0.0377807
R6430 dvdd.n520 dvdd 0.0377807
R6431 dvdd.n519 dvdd 0.0377807
R6432 dvdd.n516 dvdd 0.0377807
R6433 dvdd.n256 dvdd 0.0226354
R6434 dvdd dvdd.n266 0.0226354
R6435 dvdd.n117 dvdd 0.0226354
R6436 dvdd dvdd.n127 0.0226354
R6437 dvdd.n173 dvdd 0.0226354
R6438 dvdd dvdd.n183 0.0226354
R6439 dvdd.n331 dvdd 0.0226354
R6440 dvdd.n340 dvdd 0.0226354
R6441 dvdd dvdd.n350 0.0226354
R6442 osc_ck.n1 osc_ck.t2 236.361
R6443 osc_ck.n4 osc_ck.n2 214.567
R6444 osc_ck.n1 osc_ck.n0 207.792
R6445 osc_ck.n5 osc_ck.t0 88.3503
R6446 osc_ck.n4 osc_ck.n3 70.9231
R6447 osc_ck.n2 osc_ck.t4 29.5505
R6448 osc_ck.n2 osc_ck.t3 29.5505
R6449 osc_ck.n0 osc_ck.t1 28.5655
R6450 osc_ck.n0 osc_ck.t6 28.5655
R6451 osc_ck.n3 osc_ck.t7 18.0005
R6452 osc_ck.n3 osc_ck.t5 18.0005
R6453 osc_ck osc_ck.n5 9.94118
R6454 osc_ck.n5 osc_ck.n4 7.92796
R6455 osc_ck osc_ck.n1 3.48967
R6456 dvss.n1215 dvss.n1071 198880
R6457 dvss.n910 dvss.n909 198880
R6458 dvss.t377 dvss.n909 192115
R6459 dvss.n1215 dvss.t273 192115
R6460 dvss.n4033 dvss.n4032 82533.9
R6461 dvss.n4030 dvss.n4008 75132.3
R6462 dvss.n4009 dvss.n4008 75132.3
R6463 dvss.n4030 dvss.n4014 75132.3
R6464 dvss.n4014 dvss.n4009 75132.3
R6465 dvss.n2320 dvss.n352 48501.6
R6466 dvss.n1232 dvss.n1231 37048
R6467 dvss.n912 dvss.n911 36865.5
R6468 dvss.n4011 dvss.n3993 12828.2
R6469 dvss.n4034 dvss.n3993 12828.2
R6470 dvss.n4011 dvss.n4007 12822.4
R6471 dvss.n4034 dvss.n4007 12822.4
R6472 dvss.n235 dvss 12161.8
R6473 dvss.n176 dvss.n175 9438.11
R6474 dvss.n4054 dvss.n307 8941.81
R6475 dvss.n61 dvss.n41 8034.33
R6476 dvss.n3931 dvss.t8 8003.11
R6477 dvss.n3896 dvss.t367 8003.11
R6478 dvss.t329 dvss.n2987 8003.11
R6479 dvss.t60 dvss.n600 8003.11
R6480 dvss.t437 dvss.n2158 8003.11
R6481 dvss.n1898 dvss.t311 8003.11
R6482 dvss.t650 dvss.n1609 8003.11
R6483 dvss.n1423 dvss.t351 8003.11
R6484 dvss.t151 dvss.n1124 8003.11
R6485 dvss.t4 dvss.t2 7626.67
R6486 dvss.t6 dvss.t8 7626.67
R6487 dvss.t363 dvss.t361 7626.67
R6488 dvss.t365 dvss.t367 7626.67
R6489 dvss.t325 dvss.t323 7626.67
R6490 dvss.t329 dvss.t327 7626.67
R6491 dvss.t56 dvss.t54 7626.67
R6492 dvss.t60 dvss.t58 7626.67
R6493 dvss.t441 dvss.t445 7626.67
R6494 dvss.t437 dvss.t439 7626.67
R6495 dvss.t313 dvss.t315 7626.67
R6496 dvss.t319 dvss.t311 7626.67
R6497 dvss.t644 dvss.t646 7626.67
R6498 dvss.t650 dvss.t642 7626.67
R6499 dvss.t347 dvss.t345 7626.67
R6500 dvss.t353 dvss.t351 7626.67
R6501 dvss.t153 dvss.t149 7626.67
R6502 dvss.t151 dvss.t157 7626.67
R6503 dvss.n3721 dvss.n3720 6332.05
R6504 dvss.n3637 dvss.n498 6332.05
R6505 dvss.n2201 dvss.n2136 6332.05
R6506 dvss.n2176 dvss.n2142 6332.05
R6507 dvss.n2148 dvss.n2147 6332.05
R6508 dvss.n1979 dvss.n734 6332.05
R6509 dvss.n1599 dvss.n1598 6332.05
R6510 dvss.n1504 dvss.n843 6332.05
R6511 dvss.n1675 dvss.t200 6153.5
R6512 dvss.n3153 dvss.t200 6153.5
R6513 dvss.n3970 dvss.t663 6153.5
R6514 dvss.n3810 dvss.t180 6153.5
R6515 dvss.t200 dvss.n638 6153.5
R6516 dvss.n1966 dvss.t200 6153.5
R6517 dvss.n1491 dvss.t200 6153.5
R6518 dvss.n178 dvss.n60 5792.85
R6519 dvss.n4056 dvss.n4055 5772.37
R6520 dvss.n4055 dvss.n4054 5605.26
R6521 dvss.n235 dvss.n41 5502.51
R6522 dvss.n3970 dvss.n329 5082
R6523 dvss.n3810 dvss.n3809 5082
R6524 dvss.n3624 dvss.n508 5082
R6525 dvss.n3625 dvss.n3624 5082
R6526 dvss.n2934 dvss.n576 5082
R6527 dvss.n2198 dvss.n576 5082
R6528 dvss.n2173 dvss.n638 5082
R6529 dvss.n3153 dvss.n3152 5082
R6530 dvss.n1967 dvss.n1966 5082
R6531 dvss.n1675 dvss.n1674 5082
R6532 dvss.n1492 dvss.n1491 5082
R6533 dvss.n4029 dvss.n4015 4881.69
R6534 dvss.n4027 dvss.n4015 4881.69
R6535 dvss.n4029 dvss.n4028 4881.69
R6536 dvss.n4028 dvss.n4027 4881.69
R6537 dvss.n178 dvss.n177 4826.37
R6538 dvss.t624 dvss.n179 4465.22
R6539 dvss.n910 dvss.t379 4455
R6540 dvss.t275 dvss.n1071 4455
R6541 dvss.n59 dvss.n42 4160.18
R6542 dvss.n55 dvss.n42 4160.18
R6543 dvss.n59 dvss.n43 4160.18
R6544 dvss.n55 dvss.n43 4160.18
R6545 dvss.n175 dvss.n61 3708.43
R6546 dvss.n179 dvss.n178 3328.76
R6547 dvss.n177 dvss.n176 2962.09
R6548 dvss dvss.n61 2800
R6549 dvss.n175 dvss 2763.24
R6550 dvss.t379 dvss.t377 2310
R6551 dvss.t273 dvss.t275 2310
R6552 dvss.t374 dvss.n906 2079.65
R6553 dvss.n4033 dvss.t384 2014.07
R6554 dvss.n179 dvss.t90 1808.05
R6555 dvss.t665 dvss.t659 1778.24
R6556 dvss.t182 dvss.t174 1778.24
R6557 dvss dvss.t515 1681.61
R6558 dvss.n3931 dvss.t665 1652.85
R6559 dvss.t174 dvss.n3896 1652.85
R6560 dvss.n4012 dvss.t145 1589.55
R6561 dvss.n177 dvss.t707 1395.12
R6562 dvss.n176 dvss.t410 1376.81
R6563 dvss dvss.t162 1297.56
R6564 dvss.t453 dvss 1280.53
R6565 dvss.n54 dvss.n41 1258.81
R6566 dvss.n60 dvss.t94 1124.77
R6567 dvss.n54 dvss.t218 1124.77
R6568 dvss.t90 dvss.t70 1062.07
R6569 dvss.t70 dvss.t92 1062.07
R6570 dvss.t92 dvss.t72 1062.07
R6571 dvss.t72 dvss.t84 1062.07
R6572 dvss.t84 dvss.t76 1062.07
R6573 dvss.t76 dvss.t78 1062.07
R6574 dvss.t78 dvss.t66 1062.07
R6575 dvss.t66 dvss.t88 1062.07
R6576 dvss.t88 dvss.t62 1062.07
R6577 dvss.t62 dvss.t80 1062.07
R6578 dvss.t64 dvss.t82 1062.07
R6579 dvss.t82 dvss.t74 1062.07
R6580 dvss.t74 dvss.t86 1062.07
R6581 dvss.t86 dvss.t68 1062.07
R6582 dvss.t515 dvss.t305 1062.07
R6583 dvss.t305 dvss.t517 1062.07
R6584 dvss.t517 dvss.t303 1062.07
R6585 dvss.t68 dvss 986.207
R6586 dvss.t303 dvss 948.277
R6587 dvss.t691 dvss.t94 920.795
R6588 dvss.t307 dvss.t691 920.795
R6589 dvss.t220 dvss.t307 920.795
R6590 dvss.t218 dvss.t220 920.795
R6591 dvss.t374 dvss.n907 867.946
R6592 dvss.t235 dvss.n908 867.946
R6593 dvss dvss.n235 847.126
R6594 dvss.n4036 dvss.n4035 833.506
R6595 dvss.n4036 dvss.n3992 833.506
R6596 dvss.n4035 dvss.n4006 833.13
R6597 dvss.n4006 dvss.n3992 833.13
R6598 dvss.t719 dvss.t707 819.513
R6599 dvss.t709 dvss.t719 819.513
R6600 dvss.t721 dvss.t709 819.513
R6601 dvss.t701 dvss.t721 819.513
R6602 dvss.t725 dvss.t701 819.513
R6603 dvss.t727 dvss.t725 819.513
R6604 dvss.t715 dvss.t727 819.513
R6605 dvss.t705 dvss.t715 819.513
R6606 dvss.t711 dvss.t705 819.513
R6607 dvss.t729 dvss.t711 819.513
R6608 dvss.t713 dvss.t699 819.513
R6609 dvss.t699 dvss.t723 819.513
R6610 dvss.t723 dvss.t703 819.513
R6611 dvss.t703 dvss.t717 819.513
R6612 dvss.t162 dvss.t164 819.513
R6613 dvss.t164 dvss.t160 819.513
R6614 dvss.t160 dvss.t166 819.513
R6615 dvss.t390 dvss.t410 808.754
R6616 dvss.t412 dvss.t390 808.754
R6617 dvss.t392 dvss.t412 808.754
R6618 dvss.t404 dvss.t392 808.754
R6619 dvss.t396 dvss.t404 808.754
R6620 dvss.t398 dvss.t396 808.754
R6621 dvss.t386 dvss.t398 808.754
R6622 dvss.t408 dvss.t386 808.754
R6623 dvss.t414 dvss.t408 808.754
R6624 dvss.t400 dvss.t414 808.754
R6625 dvss.t402 dvss.t416 808.754
R6626 dvss.t394 dvss.t402 808.754
R6627 dvss.t406 dvss.t394 808.754
R6628 dvss.t388 dvss.t406 808.754
R6629 dvss.t451 dvss.t453 808.754
R6630 dvss.t447 dvss.t451 808.754
R6631 dvss.t449 dvss.t447 808.754
R6632 dvss.n4047 dvss.n307 769.572
R6633 dvss.n964 dvss.n963 769.572
R6634 dvss.n1056 dvss.n1055 769.572
R6635 dvss.n3931 dvss.t143 761.905
R6636 dvss.n3896 dvss.t477 761.905
R6637 dvss.n2987 dvss.t194 761.905
R6638 dvss.t24 dvss.n600 761.905
R6639 dvss.n2158 dvss.t630 761.905
R6640 dvss.n1898 dvss.t456 761.905
R6641 dvss.n1609 dvss.t671 761.905
R6642 dvss.n1423 dvss.t503 761.905
R6643 dvss.n1124 dvss.t422 761.905
R6644 dvss.t717 dvss 760.976
R6645 dvss dvss.t388 750.986
R6646 dvss.n3816 dvss.n428 747.437
R6647 dvss.n3561 dvss.n3560 747.437
R6648 dvss.n3409 dvss.n573 747.437
R6649 dvss.n3306 dvss.n631 747.437
R6650 dvss.n3186 dvss.n688 747.437
R6651 dvss.n1873 dvss.n1861 747.437
R6652 dvss.n1708 dvss.n797 747.437
R6653 dvss.n1398 dvss.n1386 747.437
R6654 dvss.t233 dvss.t235 745.433
R6655 dvss.t166 dvss 731.707
R6656 dvss dvss.t449 722.101
R6657 dvss.n236 dvss.t64 682.76
R6658 dvss.n909 dvss.t501 610.777
R6659 dvss.n3900 dvss.n3899 607.51
R6660 dvss.n3924 dvss.n299 607.51
R6661 dvss.n3897 dvss.t182 604.145
R6662 dvss.n3898 dvss.n350 592.001
R6663 dvss.n3925 dvss.n298 592.001
R6664 dvss.n3726 dvss.n3725 590.068
R6665 dvss.n3651 dvss.n3650 590.068
R6666 dvss.n2205 dvss.n2204 590.068
R6667 dvss.n2180 dvss.n2179 590.068
R6668 dvss.n2153 dvss.n2152 590.068
R6669 dvss.n1993 dvss.n1992 590.068
R6670 dvss.n1604 dvss.n1603 590.068
R6671 dvss.n1518 dvss.n1517 590.068
R6672 dvss.n1115 dvss.n1108 590.068
R6673 dvss.n3926 dvss.n3923 588.516
R6674 dvss.n3729 dvss.n3716 587.271
R6675 dvss.n3664 dvss.n489 587.271
R6676 dvss.n2208 dvss.n2131 587.271
R6677 dvss.n2183 dvss.n2137 587.271
R6678 dvss.n2156 dvss.n2143 587.271
R6679 dvss.n2006 dvss.n725 587.271
R6680 dvss.n1607 dvss.n1594 587.271
R6681 dvss.n1531 dvss.n834 587.271
R6682 dvss.n1182 dvss.n1181 587.271
R6683 dvss.n1514 dvss.n1513 585
R6684 dvss.n1515 dvss.n1514 585
R6685 dvss.n842 dvss.n841 585
R6686 dvss.n1516 dvss.n842 585
R6687 dvss.n1519 dvss.n1518 585
R6688 dvss.n837 dvss.n836 585
R6689 dvss.n836 dvss.n835 585
R6690 dvss.n1529 dvss.n1528 585
R6691 dvss.n1530 dvss.n1529 585
R6692 dvss.n834 dvss.n833 585
R6693 dvss.n1535 dvss.n1534 585
R6694 dvss.n1534 dvss.n1533 585
R6695 dvss.n827 dvss.n826 585
R6696 dvss.n1532 dvss.n826 585
R6697 dvss.n1544 dvss.n1543 585
R6698 dvss.n1545 dvss.n1544 585
R6699 dvss.n825 dvss.n824 585
R6700 dvss.n1546 dvss.n825 585
R6701 dvss.n1550 dvss.n1549 585
R6702 dvss.n1549 dvss.n1548 585
R6703 dvss.n819 dvss.n818 585
R6704 dvss.n1547 dvss.n818 585
R6705 dvss.n1559 dvss.n1558 585
R6706 dvss.n1560 dvss.n1559 585
R6707 dvss.n817 dvss.n816 585
R6708 dvss.n1561 dvss.n817 585
R6709 dvss.n1564 dvss.n1563 585
R6710 dvss.n1563 dvss.n1562 585
R6711 dvss.n814 dvss.n812 585
R6712 dvss.n812 dvss.n810 585
R6713 dvss.n1672 dvss.n1671 585
R6714 dvss.n1673 dvss.n1672 585
R6715 dvss.n815 dvss.n813 585
R6716 dvss.n813 dvss.n811 585
R6717 dvss.n1667 dvss.n1567 585
R6718 dvss.n1666 dvss.n1568 585
R6719 dvss.n1595 dvss.n1569 585
R6720 dvss.n1662 dvss.n1570 585
R6721 dvss.n1661 dvss.n1571 585
R6722 dvss.n1600 dvss.n1571 585
R6723 dvss.n1602 dvss.n1572 585
R6724 dvss.n1602 dvss.n1601 585
R6725 dvss.n1603 dvss.n1575 585
R6726 dvss.n1653 dvss.n1576 585
R6727 dvss.n1605 dvss.n1576 585
R6728 dvss.n1652 dvss.n1577 585
R6729 dvss.n1606 dvss.n1577 585
R6730 dvss.n1594 dvss.n1578 585
R6731 dvss.n1644 dvss.n1582 585
R6732 dvss.n1610 dvss.n1582 585
R6733 dvss.n1643 dvss.n1583 585
R6734 dvss.n1611 dvss.n1583 585
R6735 dvss.n1612 dvss.n1584 585
R6736 dvss.n1613 dvss.n1612 585
R6737 dvss.n1636 dvss.n1586 585
R6738 dvss.n1614 dvss.n1586 585
R6739 dvss.n1635 dvss.n1587 585
R6740 dvss.n1615 dvss.n1587 585
R6741 dvss.n1617 dvss.n1588 585
R6742 dvss.n1617 dvss.n1616 585
R6743 dvss.n1618 dvss.n1592 585
R6744 dvss.n1619 dvss.n1618 585
R6745 dvss.n1626 dvss.n1593 585
R6746 dvss.n1620 dvss.n1593 585
R6747 dvss.n1625 dvss.n1622 585
R6748 dvss.n1622 dvss.n1621 585
R6749 dvss.n742 dvss.n741 585
R6750 dvss.n743 dvss.n742 585
R6751 dvss.n1971 dvss.n1970 585
R6752 dvss.n1970 dvss.n1969 585
R6753 dvss.n740 dvss.n739 585
R6754 dvss.n1968 dvss.n739 585
R6755 dvss.n1977 dvss.n1976 585
R6756 dvss.n738 dvss.n737 585
R6757 dvss.n1982 dvss.n1981 585
R6758 dvss.n736 dvss.n735 585
R6759 dvss.n1989 dvss.n1988 585
R6760 dvss.n1990 dvss.n1989 585
R6761 dvss.n733 dvss.n732 585
R6762 dvss.n1991 dvss.n733 585
R6763 dvss.n1994 dvss.n1993 585
R6764 dvss.n728 dvss.n727 585
R6765 dvss.n727 dvss.n726 585
R6766 dvss.n2004 dvss.n2003 585
R6767 dvss.n2005 dvss.n2004 585
R6768 dvss.n725 dvss.n724 585
R6769 dvss.n2010 dvss.n2009 585
R6770 dvss.n2009 dvss.n2008 585
R6771 dvss.n718 dvss.n717 585
R6772 dvss.n2007 dvss.n717 585
R6773 dvss.n2019 dvss.n2018 585
R6774 dvss.n2020 dvss.n2019 585
R6775 dvss.n716 dvss.n715 585
R6776 dvss.n2021 dvss.n716 585
R6777 dvss.n2025 dvss.n2024 585
R6778 dvss.n2024 dvss.n2023 585
R6779 dvss.n710 dvss.n709 585
R6780 dvss.n2022 dvss.n709 585
R6781 dvss.n2034 dvss.n2033 585
R6782 dvss.n2035 dvss.n2034 585
R6783 dvss.n708 dvss.n707 585
R6784 dvss.n2036 dvss.n708 585
R6785 dvss.n2039 dvss.n2038 585
R6786 dvss.n2038 dvss.n2037 585
R6787 dvss.n705 dvss.n703 585
R6788 dvss.n703 dvss.n701 585
R6789 dvss.n3150 dvss.n3149 585
R6790 dvss.n3151 dvss.n3150 585
R6791 dvss.n706 dvss.n704 585
R6792 dvss.n704 dvss.n702 585
R6793 dvss.n3145 dvss.n2042 585
R6794 dvss.n3144 dvss.n2043 585
R6795 dvss.n2144 dvss.n2044 585
R6796 dvss.n3140 dvss.n2045 585
R6797 dvss.n3139 dvss.n2046 585
R6798 dvss.n2149 dvss.n2046 585
R6799 dvss.n2151 dvss.n2047 585
R6800 dvss.n2151 dvss.n2150 585
R6801 dvss.n2152 dvss.n2050 585
R6802 dvss.n3131 dvss.n2051 585
R6803 dvss.n2154 dvss.n2051 585
R6804 dvss.n3130 dvss.n2052 585
R6805 dvss.n2155 dvss.n2052 585
R6806 dvss.n2143 dvss.n2053 585
R6807 dvss.n3122 dvss.n2057 585
R6808 dvss.n2159 dvss.n2057 585
R6809 dvss.n3121 dvss.n2058 585
R6810 dvss.n2160 dvss.n2058 585
R6811 dvss.n2161 dvss.n2059 585
R6812 dvss.n2162 dvss.n2161 585
R6813 dvss.n3114 dvss.n2061 585
R6814 dvss.n2163 dvss.n2061 585
R6815 dvss.n3113 dvss.n2062 585
R6816 dvss.n2164 dvss.n2062 585
R6817 dvss.n2166 dvss.n2063 585
R6818 dvss.n2166 dvss.n2165 585
R6819 dvss.n2167 dvss.n2067 585
R6820 dvss.n2168 dvss.n2167 585
R6821 dvss.n3104 dvss.n2068 585
R6822 dvss.n2169 dvss.n2068 585
R6823 dvss.n3103 dvss.n2069 585
R6824 dvss.n2170 dvss.n2069 585
R6825 dvss.n2171 dvss.n2070 585
R6826 dvss.n2172 dvss.n2171 585
R6827 dvss.n3099 dvss.n2071 585
R6828 dvss.n2174 dvss.n2071 585
R6829 dvss.n3098 dvss.n2072 585
R6830 dvss.n2175 dvss.n2072 585
R6831 dvss.n2140 dvss.n2073 585
R6832 dvss.n3094 dvss.n2074 585
R6833 dvss.n3093 dvss.n2075 585
R6834 dvss.n2138 dvss.n2076 585
R6835 dvss.n3089 dvss.n2077 585
R6836 dvss.n2177 dvss.n2077 585
R6837 dvss.n3088 dvss.n2078 585
R6838 dvss.n2178 dvss.n2078 585
R6839 dvss.n2179 dvss.n2079 585
R6840 dvss.n3081 dvss.n2082 585
R6841 dvss.n2181 dvss.n2082 585
R6842 dvss.n3080 dvss.n2083 585
R6843 dvss.n2182 dvss.n2083 585
R6844 dvss.n2137 dvss.n2084 585
R6845 dvss.n3072 dvss.n2088 585
R6846 dvss.n2184 dvss.n2088 585
R6847 dvss.n3071 dvss.n2089 585
R6848 dvss.n2185 dvss.n2089 585
R6849 dvss.n2186 dvss.n2090 585
R6850 dvss.n2187 dvss.n2186 585
R6851 dvss.n3064 dvss.n2092 585
R6852 dvss.n2188 dvss.n2092 585
R6853 dvss.n3063 dvss.n2093 585
R6854 dvss.n2189 dvss.n2093 585
R6855 dvss.n2191 dvss.n2094 585
R6856 dvss.n2191 dvss.n2190 585
R6857 dvss.n2192 dvss.n2098 585
R6858 dvss.n2193 dvss.n2192 585
R6859 dvss.n3054 dvss.n2099 585
R6860 dvss.n2194 dvss.n2099 585
R6861 dvss.n3053 dvss.n2100 585
R6862 dvss.n2195 dvss.n2100 585
R6863 dvss.n2196 dvss.n2101 585
R6864 dvss.n2197 dvss.n2196 585
R6865 dvss.n3049 dvss.n2102 585
R6866 dvss.n2199 dvss.n2102 585
R6867 dvss.n3048 dvss.n2103 585
R6868 dvss.n2200 dvss.n2103 585
R6869 dvss.n2134 dvss.n2104 585
R6870 dvss.n3044 dvss.n2105 585
R6871 dvss.n3043 dvss.n2106 585
R6872 dvss.n2132 dvss.n2107 585
R6873 dvss.n3039 dvss.n2108 585
R6874 dvss.n2202 dvss.n2108 585
R6875 dvss.n3038 dvss.n2109 585
R6876 dvss.n2203 dvss.n2109 585
R6877 dvss.n2204 dvss.n2110 585
R6878 dvss.n3031 dvss.n2113 585
R6879 dvss.n2206 dvss.n2113 585
R6880 dvss.n3030 dvss.n2114 585
R6881 dvss.n2207 dvss.n2114 585
R6882 dvss.n2131 dvss.n2115 585
R6883 dvss.n3022 dvss.n2119 585
R6884 dvss.n2988 dvss.n2119 585
R6885 dvss.n3021 dvss.n2120 585
R6886 dvss.n2989 dvss.n2120 585
R6887 dvss.n2990 dvss.n2121 585
R6888 dvss.n2991 dvss.n2990 585
R6889 dvss.n3014 dvss.n2123 585
R6890 dvss.n2992 dvss.n2123 585
R6891 dvss.n3013 dvss.n2124 585
R6892 dvss.n2993 dvss.n2124 585
R6893 dvss.n2995 dvss.n2125 585
R6894 dvss.n2995 dvss.n2994 585
R6895 dvss.n2996 dvss.n2129 585
R6896 dvss.n2997 dvss.n2996 585
R6897 dvss.n3004 dvss.n2130 585
R6898 dvss.n2998 dvss.n2130 585
R6899 dvss.n3003 dvss.n3000 585
R6900 dvss.n3000 dvss.n2999 585
R6901 dvss.n506 dvss.n505 585
R6902 dvss.n507 dvss.n506 585
R6903 dvss.n3629 dvss.n3628 585
R6904 dvss.n3628 dvss.n3627 585
R6905 dvss.n504 dvss.n503 585
R6906 dvss.n3626 dvss.n503 585
R6907 dvss.n3635 dvss.n3634 585
R6908 dvss.n502 dvss.n501 585
R6909 dvss.n3640 dvss.n3639 585
R6910 dvss.n500 dvss.n499 585
R6911 dvss.n3647 dvss.n3646 585
R6912 dvss.n3648 dvss.n3647 585
R6913 dvss.n497 dvss.n496 585
R6914 dvss.n3649 dvss.n497 585
R6915 dvss.n3652 dvss.n3651 585
R6916 dvss.n492 dvss.n491 585
R6917 dvss.n491 dvss.n490 585
R6918 dvss.n3662 dvss.n3661 585
R6919 dvss.n3663 dvss.n3662 585
R6920 dvss.n489 dvss.n488 585
R6921 dvss.n3668 dvss.n3667 585
R6922 dvss.n3667 dvss.n3666 585
R6923 dvss.n482 dvss.n481 585
R6924 dvss.n3665 dvss.n481 585
R6925 dvss.n3677 dvss.n3676 585
R6926 dvss.n3678 dvss.n3677 585
R6927 dvss.n480 dvss.n479 585
R6928 dvss.n3679 dvss.n480 585
R6929 dvss.n3683 dvss.n3682 585
R6930 dvss.n3682 dvss.n3681 585
R6931 dvss.n474 dvss.n473 585
R6932 dvss.n3680 dvss.n473 585
R6933 dvss.n3692 dvss.n3691 585
R6934 dvss.n3693 dvss.n3692 585
R6935 dvss.n472 dvss.n471 585
R6936 dvss.n3694 dvss.n472 585
R6937 dvss.n3697 dvss.n3696 585
R6938 dvss.n3696 dvss.n3695 585
R6939 dvss.n469 dvss.n467 585
R6940 dvss.n467 dvss.n465 585
R6941 dvss.n3807 dvss.n3806 585
R6942 dvss.n3808 dvss.n3807 585
R6943 dvss.n470 dvss.n468 585
R6944 dvss.n468 dvss.n466 585
R6945 dvss.n3802 dvss.n3700 585
R6946 dvss.n3801 dvss.n3701 585
R6947 dvss.n3717 dvss.n3702 585
R6948 dvss.n3797 dvss.n3703 585
R6949 dvss.n3796 dvss.n3704 585
R6950 dvss.n3722 dvss.n3704 585
R6951 dvss.n3724 dvss.n3705 585
R6952 dvss.n3724 dvss.n3723 585
R6953 dvss.n3725 dvss.n3708 585
R6954 dvss.n3788 dvss.n3709 585
R6955 dvss.n3727 dvss.n3709 585
R6956 dvss.n3787 dvss.n3710 585
R6957 dvss.n3728 dvss.n3710 585
R6958 dvss.n3716 dvss.n3711 585
R6959 dvss.n3779 dvss.n3715 585
R6960 dvss.n3730 dvss.n3715 585
R6961 dvss.n3778 dvss.n3732 585
R6962 dvss.n3732 dvss.n3731 585
R6963 dvss.n3744 dvss.n3733 585
R6964 dvss.n3745 dvss.n3744 585
R6965 dvss.n3771 dvss.n3735 585
R6966 dvss.n3746 dvss.n3735 585
R6967 dvss.n3770 dvss.n3736 585
R6968 dvss.n3747 dvss.n3736 585
R6969 dvss.n3749 dvss.n3737 585
R6970 dvss.n3749 dvss.n3748 585
R6971 dvss.n3750 dvss.n3741 585
R6972 dvss.n3751 dvss.n3750 585
R6973 dvss.n3761 dvss.n3742 585
R6974 dvss.n3752 dvss.n3742 585
R6975 dvss.n3760 dvss.n3743 585
R6976 dvss.n3753 dvss.n3743 585
R6977 dvss.n3756 dvss.n3755 585
R6978 dvss.n3755 dvss.n3754 585
R6979 dvss.n311 dvss.n309 585
R6980 dvss.n309 dvss.n308 585
R6981 dvss.n4052 dvss.n4051 585
R6982 dvss.n4053 dvss.n4052 585
R6983 dvss.n312 dvss.n310 585
R6984 dvss.n1502 dvss.n1501 585
R6985 dvss.n847 dvss.n846 585
R6986 dvss.n1507 dvss.n1506 585
R6987 dvss.n845 dvss.n844 585
R6988 dvss.n1107 dvss.n1106 585
R6989 dvss.n1191 dvss.n1107 585
R6990 dvss.n1189 dvss.n1188 585
R6991 dvss.n1190 dvss.n1189 585
R6992 dvss.n1187 dvss.n1108 585
R6993 dvss.n1186 dvss.n1185 585
R6994 dvss.n1185 dvss.n1184 585
R6995 dvss.n1114 dvss.n1113 585
R6996 dvss.n1183 dvss.n1114 585
R6997 dvss.n1181 dvss.n1180 585
R6998 dvss.n1179 dvss.n1116 585
R6999 dvss.n1122 dvss.n1116 585
R7000 dvss.n1178 dvss.n1177 585
R7001 dvss.n1177 dvss.n1176 585
R7002 dvss.n1121 dvss.n1120 585
R7003 dvss.n1175 dvss.n1121 585
R7004 dvss.n1173 dvss.n1172 585
R7005 dvss.n1174 dvss.n1173 585
R7006 dvss.n1171 dvss.n1126 585
R7007 dvss.n1126 dvss.n1125 585
R7008 dvss.n1170 dvss.n1169 585
R7009 dvss.n1169 dvss.n1168 585
R7010 dvss.n1149 dvss.n1148 585
R7011 dvss.n1167 dvss.n1149 585
R7012 dvss.n1165 dvss.n1164 585
R7013 dvss.n1166 dvss.n1165 585
R7014 dvss.n1163 dvss.n1151 585
R7015 dvss.n1151 dvss.n1150 585
R7016 dvss.n851 dvss.n850 585
R7017 dvss.n852 dvss.n851 585
R7018 dvss.n1496 dvss.n1495 585
R7019 dvss.n1495 dvss.n1494 585
R7020 dvss.n849 dvss.n848 585
R7021 dvss.n1493 dvss.n848 585
R7022 dvss.n900 dvss.n899 585
R7023 dvss.n1234 dvss.n899 585
R7024 dvss.n1246 dvss.n1245 585
R7025 dvss.n1247 dvss.n1246 585
R7026 dvss.n896 dvss.n895 585
R7027 dvss.n1248 dvss.n895 585
R7028 dvss.n1259 dvss.n1258 585
R7029 dvss.n1259 dvss.n893 585
R7030 dvss.n1260 dvss.n888 585
R7031 dvss.n1261 dvss.n1260 585
R7032 dvss.n1273 dvss.n889 585
R7033 dvss.n894 dvss.n889 585
R7034 dvss.n1274 dvss.n884 585
R7035 dvss.n1279 dvss.n884 585
R7036 dvss.n1283 dvss.n885 585
R7037 dvss.n1283 dvss.n1282 585
R7038 dvss.n1284 dvss.n879 585
R7039 dvss.n1285 dvss.n1284 585
R7040 dvss.n1294 dvss.n880 585
R7041 dvss.n1123 dvss.n880 585
R7042 dvss.n1295 dvss.n874 585
R7043 dvss.n876 dvss.n874 585
R7044 dvss.n1308 dvss.n875 585
R7045 dvss.n1308 dvss.n1307 585
R7046 dvss.n1309 dvss.n867 585
R7047 dvss.n1310 dvss.n1309 585
R7048 dvss.n873 dvss.n872 585
R7049 dvss.n1311 dvss.n873 585
R7050 dvss.n1315 dvss.n1314 585
R7051 dvss.n1314 dvss.n1313 585
R7052 dvss.n858 dvss.n856 585
R7053 dvss.n856 dvss.n853 585
R7054 dvss.n1489 dvss.n1488 585
R7055 dvss.n1490 dvss.n1489 585
R7056 dvss.n859 dvss.n857 585
R7057 dvss.n857 dvss.n855 585
R7058 dvss.n1396 dvss.n1330 585
R7059 dvss.n1395 dvss.n1331 585
R7060 dvss.n1394 dvss.n1335 585
R7061 dvss.n1400 dvss.n1336 585
R7062 dvss.n1402 dvss.n1401 585
R7063 dvss.n1403 dvss.n1402 585
R7064 dvss.n1385 dvss.n1340 585
R7065 dvss.n1404 dvss.n1385 585
R7066 dvss.n1406 dvss.n1345 585
R7067 dvss.n1406 dvss.n1405 585
R7068 dvss.n1408 dvss.n1407 585
R7069 dvss.n1407 dvss.n1382 585
R7070 dvss.n1412 dvss.n1411 585
R7071 dvss.n1413 dvss.n1412 585
R7072 dvss.n1381 dvss.n1351 585
R7073 dvss.n1414 dvss.n1381 585
R7074 dvss.n1417 dvss.n1356 585
R7075 dvss.n1417 dvss.n1416 585
R7076 dvss.n1418 dvss.n1357 585
R7077 dvss.n1419 dvss.n1418 585
R7078 dvss.n1379 dvss.n1378 585
R7079 dvss.n1422 dvss.n1379 585
R7080 dvss.n1425 dvss.n1360 585
R7081 dvss.n1425 dvss.n1424 585
R7082 dvss.n1426 dvss.n1368 585
R7083 dvss.n1427 dvss.n1426 585
R7084 dvss.n1376 dvss.n1369 585
R7085 dvss.n1428 dvss.n1376 585
R7086 dvss.n1432 dvss.n1377 585
R7087 dvss.n1432 dvss.n1431 585
R7088 dvss.n1433 dvss.n1373 585
R7089 dvss.n1434 dvss.n1433 585
R7090 dvss.n808 dvss.n807 585
R7091 dvss.n1435 dvss.n808 585
R7092 dvss.n1678 dvss.n1677 585
R7093 dvss.n1677 dvss.n1676 585
R7094 dvss.n802 dvss.n800 585
R7095 dvss.n800 dvss.n798 585
R7096 dvss.n1706 dvss.n1705 585
R7097 dvss.n1707 dvss.n1706 585
R7098 dvss.n803 dvss.n801 585
R7099 dvss.n1694 dvss.n1692 585
R7100 dvss.n1698 dvss.n1697 585
R7101 dvss.n1695 dvss.n793 585
R7102 dvss.n791 dvss.n790 585
R7103 dvss.n1709 dvss.n790 585
R7104 dvss.n1721 dvss.n1720 585
R7105 dvss.n1722 dvss.n1721 585
R7106 dvss.n787 dvss.n786 585
R7107 dvss.n1723 dvss.n786 585
R7108 dvss.n1734 dvss.n1733 585
R7109 dvss.n1734 dvss.n784 585
R7110 dvss.n1735 dvss.n779 585
R7111 dvss.n1736 dvss.n1735 585
R7112 dvss.n1748 dvss.n780 585
R7113 dvss.n785 dvss.n780 585
R7114 dvss.n1749 dvss.n775 585
R7115 dvss.n1754 dvss.n775 585
R7116 dvss.n1758 dvss.n776 585
R7117 dvss.n1758 dvss.n1757 585
R7118 dvss.n1759 dvss.n770 585
R7119 dvss.n1760 dvss.n1759 585
R7120 dvss.n1769 dvss.n771 585
R7121 dvss.n1608 dvss.n771 585
R7122 dvss.n1770 dvss.n765 585
R7123 dvss.n767 dvss.n765 585
R7124 dvss.n1783 dvss.n766 585
R7125 dvss.n1783 dvss.n1782 585
R7126 dvss.n1784 dvss.n758 585
R7127 dvss.n1785 dvss.n1784 585
R7128 dvss.n764 dvss.n763 585
R7129 dvss.n1786 dvss.n764 585
R7130 dvss.n1790 dvss.n1789 585
R7131 dvss.n1789 dvss.n1788 585
R7132 dvss.n749 dvss.n747 585
R7133 dvss.n747 dvss.n744 585
R7134 dvss.n1964 dvss.n1963 585
R7135 dvss.n1965 dvss.n1964 585
R7136 dvss.n750 dvss.n748 585
R7137 dvss.n748 dvss.n746 585
R7138 dvss.n1871 dvss.n1805 585
R7139 dvss.n1870 dvss.n1806 585
R7140 dvss.n1869 dvss.n1810 585
R7141 dvss.n1875 dvss.n1811 585
R7142 dvss.n1877 dvss.n1876 585
R7143 dvss.n1878 dvss.n1877 585
R7144 dvss.n1860 dvss.n1815 585
R7145 dvss.n1879 dvss.n1860 585
R7146 dvss.n1881 dvss.n1820 585
R7147 dvss.n1881 dvss.n1880 585
R7148 dvss.n1883 dvss.n1882 585
R7149 dvss.n1882 dvss.n1857 585
R7150 dvss.n1887 dvss.n1886 585
R7151 dvss.n1888 dvss.n1887 585
R7152 dvss.n1856 dvss.n1826 585
R7153 dvss.n1889 dvss.n1856 585
R7154 dvss.n1892 dvss.n1831 585
R7155 dvss.n1892 dvss.n1891 585
R7156 dvss.n1893 dvss.n1832 585
R7157 dvss.n1894 dvss.n1893 585
R7158 dvss.n1854 dvss.n1853 585
R7159 dvss.n1897 dvss.n1854 585
R7160 dvss.n1900 dvss.n1835 585
R7161 dvss.n1900 dvss.n1899 585
R7162 dvss.n1901 dvss.n1843 585
R7163 dvss.n1902 dvss.n1901 585
R7164 dvss.n1851 dvss.n1844 585
R7165 dvss.n1903 dvss.n1851 585
R7166 dvss.n1907 dvss.n1852 585
R7167 dvss.n1907 dvss.n1906 585
R7168 dvss.n1908 dvss.n1848 585
R7169 dvss.n1909 dvss.n1908 585
R7170 dvss.n699 dvss.n698 585
R7171 dvss.n1910 dvss.n699 585
R7172 dvss.n3156 dvss.n3155 585
R7173 dvss.n3155 dvss.n3154 585
R7174 dvss.n693 dvss.n691 585
R7175 dvss.n691 dvss.n689 585
R7176 dvss.n3184 dvss.n3183 585
R7177 dvss.n3185 dvss.n3184 585
R7178 dvss.n694 dvss.n692 585
R7179 dvss.n3172 dvss.n3170 585
R7180 dvss.n3176 dvss.n3175 585
R7181 dvss.n3173 dvss.n684 585
R7182 dvss.n682 dvss.n681 585
R7183 dvss.n3187 dvss.n681 585
R7184 dvss.n3199 dvss.n3198 585
R7185 dvss.n3200 dvss.n3199 585
R7186 dvss.n678 dvss.n677 585
R7187 dvss.n3201 dvss.n677 585
R7188 dvss.n3212 dvss.n3211 585
R7189 dvss.n3212 dvss.n675 585
R7190 dvss.n3213 dvss.n670 585
R7191 dvss.n3214 dvss.n3213 585
R7192 dvss.n3226 dvss.n671 585
R7193 dvss.n676 dvss.n671 585
R7194 dvss.n3227 dvss.n666 585
R7195 dvss.n3232 dvss.n666 585
R7196 dvss.n3236 dvss.n667 585
R7197 dvss.n3236 dvss.n3235 585
R7198 dvss.n3237 dvss.n661 585
R7199 dvss.n3238 dvss.n3237 585
R7200 dvss.n3247 dvss.n662 585
R7201 dvss.n2157 dvss.n662 585
R7202 dvss.n3248 dvss.n656 585
R7203 dvss.n658 dvss.n656 585
R7204 dvss.n3261 dvss.n657 585
R7205 dvss.n3261 dvss.n3260 585
R7206 dvss.n3262 dvss.n649 585
R7207 dvss.n3263 dvss.n3262 585
R7208 dvss.n655 dvss.n654 585
R7209 dvss.n3264 dvss.n655 585
R7210 dvss.n3269 dvss.n3268 585
R7211 dvss.n3268 dvss.n3267 585
R7212 dvss.n640 dvss.n639 585
R7213 dvss.n3266 dvss.n639 585
R7214 dvss.n3285 dvss.n3284 585
R7215 dvss.n3286 dvss.n3285 585
R7216 dvss.n634 dvss.n633 585
R7217 dvss.n3287 dvss.n633 585
R7218 dvss.n3304 dvss.n3303 585
R7219 dvss.n635 dvss.n632 585
R7220 dvss.n629 dvss.n628 585
R7221 dvss.n3309 dvss.n3308 585
R7222 dvss.n623 dvss.n622 585
R7223 dvss.n630 dvss.n622 585
R7224 dvss.n3321 dvss.n3320 585
R7225 dvss.n3322 dvss.n3321 585
R7226 dvss.n619 dvss.n618 585
R7227 dvss.n3323 dvss.n619 585
R7228 dvss.n3329 dvss.n3328 585
R7229 dvss.n3328 dvss.n3327 585
R7230 dvss.n613 dvss.n612 585
R7231 dvss.n3326 dvss.n612 585
R7232 dvss.n3347 dvss.n3346 585
R7233 dvss.n3348 dvss.n3347 585
R7234 dvss.n607 dvss.n606 585
R7235 dvss.n609 dvss.n607 585
R7236 dvss.n3353 dvss.n3352 585
R7237 dvss.n3352 dvss.n3351 585
R7238 dvss.n602 dvss.n601 585
R7239 dvss.n608 dvss.n601 585
R7240 dvss.n3364 dvss.n3363 585
R7241 dvss.n3365 dvss.n3364 585
R7242 dvss.n597 dvss.n596 585
R7243 dvss.n596 dvss.n594 585
R7244 dvss.n3378 dvss.n3377 585
R7245 dvss.n3379 dvss.n3378 585
R7246 dvss.n592 dvss.n586 585
R7247 dvss.n3380 dvss.n592 585
R7248 dvss.n3386 dvss.n3385 585
R7249 dvss.n3385 dvss.n3384 585
R7250 dvss.n593 dvss.n580 585
R7251 dvss.n3383 dvss.n593 585
R7252 dvss.n3398 dvss.n581 585
R7253 dvss.n3382 dvss.n581 585
R7254 dvss.n3399 dvss.n574 585
R7255 dvss.n3404 dvss.n574 585
R7256 dvss.n3406 dvss.n575 585
R7257 dvss.n3406 dvss.n3405 585
R7258 dvss.n3407 dvss.n568 585
R7259 dvss.n570 dvss.n569 585
R7260 dvss.n3412 dvss.n3411 585
R7261 dvss.n571 dvss.n559 585
R7262 dvss.n3430 dvss.n560 585
R7263 dvss.n572 dvss.n560 585
R7264 dvss.n3431 dvss.n555 585
R7265 dvss.n3441 dvss.n555 585
R7266 dvss.n3443 dvss.n556 585
R7267 dvss.n3443 dvss.n3442 585
R7268 dvss.n3444 dvss.n550 585
R7269 dvss.n3445 dvss.n3444 585
R7270 dvss.n545 dvss.n544 585
R7271 dvss.n554 dvss.n544 585
R7272 dvss.n3463 dvss.n3462 585
R7273 dvss.n3464 dvss.n3463 585
R7274 dvss.n546 dvss.n540 585
R7275 dvss.n542 dvss.n540 585
R7276 dvss.n3468 dvss.n541 585
R7277 dvss.n3468 dvss.n3467 585
R7278 dvss.n3469 dvss.n535 585
R7279 dvss.n3470 dvss.n3469 585
R7280 dvss.n3479 dvss.n536 585
R7281 dvss.n2209 dvss.n536 585
R7282 dvss.n3480 dvss.n530 585
R7283 dvss.n532 dvss.n530 585
R7284 dvss.n3493 dvss.n531 585
R7285 dvss.n3493 dvss.n3492 585
R7286 dvss.n3494 dvss.n523 585
R7287 dvss.n3495 dvss.n3494 585
R7288 dvss.n529 dvss.n528 585
R7289 dvss.n3496 dvss.n529 585
R7290 dvss.n3500 dvss.n3499 585
R7291 dvss.n3499 dvss.n3498 585
R7292 dvss.n514 dvss.n512 585
R7293 dvss.n512 dvss.n509 585
R7294 dvss.n3622 dvss.n3621 585
R7295 dvss.n3623 dvss.n3622 585
R7296 dvss.n515 dvss.n513 585
R7297 dvss.n513 dvss.n511 585
R7298 dvss.n3558 dvss.n3515 585
R7299 dvss.n3557 dvss.n3516 585
R7300 dvss.n3556 dvss.n3520 585
R7301 dvss.n3554 dvss.n3521 585
R7302 dvss.n3553 dvss.n3552 585
R7303 dvss.n3569 dvss.n3553 585
R7304 dvss.n3571 dvss.n3525 585
R7305 dvss.n3571 dvss.n3570 585
R7306 dvss.n3572 dvss.n3530 585
R7307 dvss.n3573 dvss.n3572 585
R7308 dvss.n3548 dvss.n3547 585
R7309 dvss.n3574 dvss.n3547 585
R7310 dvss.n3578 dvss.n3551 585
R7311 dvss.n3578 dvss.n3577 585
R7312 dvss.n3579 dvss.n3536 585
R7313 dvss.n3580 dvss.n3579 585
R7314 dvss.n3542 dvss.n3541 585
R7315 dvss.n3546 dvss.n3542 585
R7316 dvss.n3585 dvss.n3584 585
R7317 dvss.n3584 dvss.n3583 585
R7318 dvss.n374 dvss.n372 585
R7319 dvss.n3543 dvss.n372 585
R7320 dvss.n3894 dvss.n3893 585
R7321 dvss.n3895 dvss.n3894 585
R7322 dvss.n375 dvss.n373 585
R7323 dvss.n445 dvss.n373 585
R7324 dvss.n444 dvss.n379 585
R7325 dvss.n446 dvss.n444 585
R7326 dvss.n452 dvss.n451 585
R7327 dvss.n451 dvss.n450 585
R7328 dvss.n455 dvss.n454 585
R7329 dvss.n456 dvss.n455 585
R7330 dvss.n441 dvss.n440 585
R7331 dvss.n457 dvss.n440 585
R7332 dvss.n463 dvss.n462 585
R7333 dvss.n464 dvss.n463 585
R7334 dvss.n438 dvss.n388 585
R7335 dvss.n3811 dvss.n438 585
R7336 dvss.n3813 dvss.n393 585
R7337 dvss.n3813 dvss.n3812 585
R7338 dvss.n3814 dvss.n394 585
R7339 dvss.n437 dvss.n395 585
R7340 dvss.n436 dvss.n399 585
R7341 dvss.n3818 dvss.n400 585
R7342 dvss.n3820 dvss.n3819 585
R7343 dvss.n3821 dvss.n3820 585
R7344 dvss.n427 dvss.n404 585
R7345 dvss.n3822 dvss.n427 585
R7346 dvss.n3824 dvss.n409 585
R7347 dvss.n3824 dvss.n3823 585
R7348 dvss.n3826 dvss.n3825 585
R7349 dvss.n3825 dvss.n424 585
R7350 dvss.n3830 dvss.n3829 585
R7351 dvss.n3831 dvss.n3830 585
R7352 dvss.n423 dvss.n415 585
R7353 dvss.n3832 dvss.n423 585
R7354 dvss.n3835 dvss.n420 585
R7355 dvss.n3835 dvss.n3834 585
R7356 dvss.n3836 dvss.n421 585
R7357 dvss.n3837 dvss.n3836 585
R7358 dvss.n349 dvss.n348 585
R7359 dvss.n3839 dvss.n349 585
R7360 dvss.n3934 dvss.n3933 585
R7361 dvss.n3933 dvss.n3932 585
R7362 dvss.n343 dvss.n342 585
R7363 dvss.n345 dvss.n343 585
R7364 dvss.n3945 dvss.n3944 585
R7365 dvss.n3944 dvss.n3943 585
R7366 dvss.n344 dvss.n338 585
R7367 dvss.n3942 dvss.n344 585
R7368 dvss.n333 dvss.n332 585
R7369 dvss.n3941 dvss.n332 585
R7370 dvss.n3965 dvss.n3964 585
R7371 dvss.n3966 dvss.n3965 585
R7372 dvss.n324 dvss.n323 585
R7373 dvss.n3969 dvss.n324 585
R7374 dvss.n3973 dvss.n3972 585
R7375 dvss.n3972 dvss.n3971 585
R7376 dvss.n319 dvss.n317 585
R7377 dvss.n317 dvss.n316 585
R7378 dvss.n3980 dvss.n3979 585
R7379 dvss.n3981 dvss.n3980 585
R7380 dvss.n318 dvss.n313 585
R7381 dvss.n318 dvss.n306 585
R7382 dvss.n1014 dvss.n935 585
R7383 dvss.n1017 dvss.n1016 585
R7384 dvss.n951 dvss.n936 585
R7385 dvss.n951 dvss.n906 585
R7386 dvss.n950 dvss.n949 585
R7387 dvss.n937 dvss.n902 585
R7388 dvss.n1030 dvss.n931 585
R7389 dvss.n943 dvss.n931 585
R7390 dvss.n941 dvss.n932 585
R7391 dvss.n946 dvss.n945 585
R7392 dvss.n940 dvss.n903 585
R7393 dvss.n1237 dvss.n904 585
R7394 dvss.n1236 dvss.n1235 585
R7395 dvss.n1235 dvss.n1234 585
R7396 dvss.n898 dvss.n897 585
R7397 dvss.n1247 dvss.n898 585
R7398 dvss.n1250 dvss.n1249 585
R7399 dvss.n1249 dvss.n1248 585
R7400 dvss.n892 dvss.n891 585
R7401 dvss.n893 dvss.n892 585
R7402 dvss.n1263 dvss.n1262 585
R7403 dvss.n1262 dvss.n1261 585
R7404 dvss.n887 dvss.n886 585
R7405 dvss.n894 dvss.n886 585
R7406 dvss.n1278 dvss.n1277 585
R7407 dvss.n1279 dvss.n1278 585
R7408 dvss.n883 dvss.n882 585
R7409 dvss.n1282 dvss.n883 585
R7410 dvss.n1287 dvss.n1286 585
R7411 dvss.n1286 dvss.n1285 585
R7412 dvss.n878 dvss.n877 585
R7413 dvss.n1123 dvss.n877 585
R7414 dvss.n1305 dvss.n1304 585
R7415 dvss.n1305 dvss.n876 585
R7416 dvss.n1306 dvss.n869 585
R7417 dvss.n1307 dvss.n1306 585
R7418 dvss.n1319 dvss.n870 585
R7419 dvss.n1310 dvss.n870 585
R7420 dvss.n1318 dvss.n871 585
R7421 dvss.n1311 dvss.n871 585
R7422 dvss.n1312 dvss.n861 585
R7423 dvss.n1313 dvss.n1312 585
R7424 dvss.n1327 dvss.n862 585
R7425 dvss.n862 dvss.n853 585
R7426 dvss.n1486 dvss.n854 585
R7427 dvss.n1490 dvss.n854 585
R7428 dvss.n1485 dvss.n1328 585
R7429 dvss.n1328 dvss.n855 585
R7430 dvss.n1388 dvss.n1329 585
R7431 dvss.n1481 dvss.n1332 585
R7432 dvss.n1480 dvss.n1333 585
R7433 dvss.n1392 dvss.n1334 585
R7434 dvss.n1393 dvss.n1341 585
R7435 dvss.n1403 dvss.n1393 585
R7436 dvss.n1473 dvss.n1342 585
R7437 dvss.n1404 dvss.n1342 585
R7438 dvss.n1472 dvss.n1343 585
R7439 dvss.n1405 dvss.n1343 585
R7440 dvss.n1383 dvss.n1344 585
R7441 dvss.n1383 dvss.n1382 585
R7442 dvss.n1384 dvss.n1352 585
R7443 dvss.n1413 dvss.n1384 585
R7444 dvss.n1464 dvss.n1353 585
R7445 dvss.n1414 dvss.n1353 585
R7446 dvss.n1463 dvss.n1354 585
R7447 dvss.n1416 dvss.n1354 585
R7448 dvss.n1420 dvss.n1355 585
R7449 dvss.n1420 dvss.n1419 585
R7450 dvss.n1421 dvss.n1361 585
R7451 dvss.n1422 dvss.n1421 585
R7452 dvss.n1453 dvss.n1362 585
R7453 dvss.n1424 dvss.n1362 585
R7454 dvss.n1452 dvss.n1363 585
R7455 dvss.n1427 dvss.n1363 585
R7456 dvss.n1429 dvss.n1364 585
R7457 dvss.n1429 dvss.n1428 585
R7458 dvss.n1430 dvss.n1374 585
R7459 dvss.n1431 dvss.n1430 585
R7460 dvss.n1439 dvss.n1375 585
R7461 dvss.n1434 dvss.n1375 585
R7462 dvss.n1438 dvss.n1436 585
R7463 dvss.n1436 dvss.n1435 585
R7464 dvss.n809 dvss.n804 585
R7465 dvss.n1676 dvss.n809 585
R7466 dvss.n1684 dvss.n805 585
R7467 dvss.n805 dvss.n798 585
R7468 dvss.n1703 dvss.n799 585
R7469 dvss.n1707 dvss.n799 585
R7470 dvss.n1702 dvss.n1685 585
R7471 dvss.n1691 dvss.n1690 585
R7472 dvss.n1686 dvss.n794 585
R7473 dvss.n1712 dvss.n795 585
R7474 dvss.n1711 dvss.n1710 585
R7475 dvss.n1710 dvss.n1709 585
R7476 dvss.n789 dvss.n788 585
R7477 dvss.n1722 dvss.n789 585
R7478 dvss.n1725 dvss.n1724 585
R7479 dvss.n1724 dvss.n1723 585
R7480 dvss.n783 dvss.n782 585
R7481 dvss.n784 dvss.n783 585
R7482 dvss.n1738 dvss.n1737 585
R7483 dvss.n1737 dvss.n1736 585
R7484 dvss.n778 dvss.n777 585
R7485 dvss.n785 dvss.n777 585
R7486 dvss.n1753 dvss.n1752 585
R7487 dvss.n1754 dvss.n1753 585
R7488 dvss.n774 dvss.n773 585
R7489 dvss.n1757 dvss.n774 585
R7490 dvss.n1762 dvss.n1761 585
R7491 dvss.n1761 dvss.n1760 585
R7492 dvss.n769 dvss.n768 585
R7493 dvss.n1608 dvss.n768 585
R7494 dvss.n1780 dvss.n1779 585
R7495 dvss.n1780 dvss.n767 585
R7496 dvss.n1781 dvss.n760 585
R7497 dvss.n1782 dvss.n1781 585
R7498 dvss.n1794 dvss.n761 585
R7499 dvss.n1785 dvss.n761 585
R7500 dvss.n1793 dvss.n762 585
R7501 dvss.n1786 dvss.n762 585
R7502 dvss.n1787 dvss.n752 585
R7503 dvss.n1788 dvss.n1787 585
R7504 dvss.n1802 dvss.n753 585
R7505 dvss.n753 dvss.n744 585
R7506 dvss.n1961 dvss.n745 585
R7507 dvss.n1965 dvss.n745 585
R7508 dvss.n1960 dvss.n1803 585
R7509 dvss.n1803 dvss.n746 585
R7510 dvss.n1863 dvss.n1804 585
R7511 dvss.n1956 dvss.n1807 585
R7512 dvss.n1955 dvss.n1808 585
R7513 dvss.n1867 dvss.n1809 585
R7514 dvss.n1868 dvss.n1816 585
R7515 dvss.n1878 dvss.n1868 585
R7516 dvss.n1948 dvss.n1817 585
R7517 dvss.n1879 dvss.n1817 585
R7518 dvss.n1947 dvss.n1818 585
R7519 dvss.n1880 dvss.n1818 585
R7520 dvss.n1858 dvss.n1819 585
R7521 dvss.n1858 dvss.n1857 585
R7522 dvss.n1859 dvss.n1827 585
R7523 dvss.n1888 dvss.n1859 585
R7524 dvss.n1939 dvss.n1828 585
R7525 dvss.n1889 dvss.n1828 585
R7526 dvss.n1938 dvss.n1829 585
R7527 dvss.n1891 dvss.n1829 585
R7528 dvss.n1895 dvss.n1830 585
R7529 dvss.n1895 dvss.n1894 585
R7530 dvss.n1896 dvss.n1836 585
R7531 dvss.n1897 dvss.n1896 585
R7532 dvss.n1928 dvss.n1837 585
R7533 dvss.n1899 dvss.n1837 585
R7534 dvss.n1927 dvss.n1838 585
R7535 dvss.n1902 dvss.n1838 585
R7536 dvss.n1904 dvss.n1839 585
R7537 dvss.n1904 dvss.n1903 585
R7538 dvss.n1905 dvss.n1849 585
R7539 dvss.n1906 dvss.n1905 585
R7540 dvss.n1914 dvss.n1850 585
R7541 dvss.n1909 dvss.n1850 585
R7542 dvss.n1913 dvss.n1911 585
R7543 dvss.n1911 dvss.n1910 585
R7544 dvss.n700 dvss.n695 585
R7545 dvss.n3154 dvss.n700 585
R7546 dvss.n3162 dvss.n696 585
R7547 dvss.n696 dvss.n689 585
R7548 dvss.n3181 dvss.n690 585
R7549 dvss.n3185 dvss.n690 585
R7550 dvss.n3180 dvss.n3163 585
R7551 dvss.n3169 dvss.n3168 585
R7552 dvss.n3164 dvss.n685 585
R7553 dvss.n3190 dvss.n686 585
R7554 dvss.n3189 dvss.n3188 585
R7555 dvss.n3188 dvss.n3187 585
R7556 dvss.n680 dvss.n679 585
R7557 dvss.n3200 dvss.n680 585
R7558 dvss.n3203 dvss.n3202 585
R7559 dvss.n3202 dvss.n3201 585
R7560 dvss.n674 dvss.n673 585
R7561 dvss.n675 dvss.n674 585
R7562 dvss.n3216 dvss.n3215 585
R7563 dvss.n3215 dvss.n3214 585
R7564 dvss.n669 dvss.n668 585
R7565 dvss.n676 dvss.n668 585
R7566 dvss.n3231 dvss.n3230 585
R7567 dvss.n3232 dvss.n3231 585
R7568 dvss.n665 dvss.n664 585
R7569 dvss.n3235 dvss.n665 585
R7570 dvss.n3240 dvss.n3239 585
R7571 dvss.n3239 dvss.n3238 585
R7572 dvss.n660 dvss.n659 585
R7573 dvss.n2157 dvss.n659 585
R7574 dvss.n3258 dvss.n3257 585
R7575 dvss.n3258 dvss.n658 585
R7576 dvss.n3259 dvss.n651 585
R7577 dvss.n3260 dvss.n3259 585
R7578 dvss.n3273 dvss.n652 585
R7579 dvss.n3263 dvss.n652 585
R7580 dvss.n3272 dvss.n653 585
R7581 dvss.n3264 dvss.n653 585
R7582 dvss.n3265 dvss.n643 585
R7583 dvss.n3267 dvss.n3265 585
R7584 dvss.n3281 dvss.n644 585
R7585 dvss.n3266 dvss.n644 585
R7586 dvss.n3282 dvss.n637 585
R7587 dvss.n3286 dvss.n637 585
R7588 dvss.n3288 dvss.n636 585
R7589 dvss.n3288 dvss.n3287 585
R7590 dvss.n3301 dvss.n3289 585
R7591 dvss.n3300 dvss.n3290 585
R7592 dvss.n3297 dvss.n3296 585
R7593 dvss.n3291 dvss.n626 585
R7594 dvss.n3317 dvss.n627 585
R7595 dvss.n630 dvss.n627 585
R7596 dvss.n3318 dvss.n620 585
R7597 dvss.n3322 dvss.n620 585
R7598 dvss.n3324 dvss.n621 585
R7599 dvss.n3324 dvss.n3323 585
R7600 dvss.n3325 dvss.n614 585
R7601 dvss.n3327 dvss.n3325 585
R7602 dvss.n3343 dvss.n615 585
R7603 dvss.n3326 dvss.n615 585
R7604 dvss.n3344 dvss.n611 585
R7605 dvss.n3348 dvss.n611 585
R7606 dvss.n610 dvss.n604 585
R7607 dvss.n610 dvss.n609 585
R7608 dvss.n3355 dvss.n605 585
R7609 dvss.n3351 dvss.n605 585
R7610 dvss.n3356 dvss.n599 585
R7611 dvss.n608 dvss.n599 585
R7612 dvss.n3366 dvss.n598 585
R7613 dvss.n3366 dvss.n3365 585
R7614 dvss.n3368 dvss.n3367 585
R7615 dvss.n3367 dvss.n594 585
R7616 dvss.n595 dvss.n588 585
R7617 dvss.n3379 dvss.n595 585
R7618 dvss.n3390 dvss.n589 585
R7619 dvss.n3380 dvss.n589 585
R7620 dvss.n3389 dvss.n590 585
R7621 dvss.n3384 dvss.n590 585
R7622 dvss.n3381 dvss.n591 585
R7623 dvss.n3383 dvss.n3381 585
R7624 dvss.n578 dvss.n577 585
R7625 dvss.n3382 dvss.n577 585
R7626 dvss.n3403 dvss.n3402 585
R7627 dvss.n3404 dvss.n3403 585
R7628 dvss.n566 dvss.n565 585
R7629 dvss.n3405 dvss.n565 585
R7630 dvss.n3417 dvss.n3416 585
R7631 dvss.n567 dvss.n564 585
R7632 dvss.n562 dvss.n561 585
R7633 dvss.n3422 dvss.n3421 585
R7634 dvss.n558 dvss.n557 585
R7635 dvss.n572 dvss.n557 585
R7636 dvss.n3440 dvss.n3439 585
R7637 dvss.n3441 dvss.n3440 585
R7638 dvss.n552 dvss.n551 585
R7639 dvss.n3442 dvss.n552 585
R7640 dvss.n3447 dvss.n3446 585
R7641 dvss.n3446 dvss.n3445 585
R7642 dvss.n553 dvss.n547 585
R7643 dvss.n554 dvss.n553 585
R7644 dvss.n3460 dvss.n543 585
R7645 dvss.n3464 dvss.n543 585
R7646 dvss.n3459 dvss.n548 585
R7647 dvss.n548 dvss.n542 585
R7648 dvss.n539 dvss.n538 585
R7649 dvss.n3467 dvss.n539 585
R7650 dvss.n3472 dvss.n3471 585
R7651 dvss.n3471 dvss.n3470 585
R7652 dvss.n534 dvss.n533 585
R7653 dvss.n2209 dvss.n533 585
R7654 dvss.n3490 dvss.n3489 585
R7655 dvss.n3490 dvss.n532 585
R7656 dvss.n3491 dvss.n525 585
R7657 dvss.n3492 dvss.n3491 585
R7658 dvss.n3504 dvss.n526 585
R7659 dvss.n3495 dvss.n526 585
R7660 dvss.n3503 dvss.n527 585
R7661 dvss.n3496 dvss.n527 585
R7662 dvss.n3497 dvss.n517 585
R7663 dvss.n3498 dvss.n3497 585
R7664 dvss.n3512 dvss.n518 585
R7665 dvss.n518 dvss.n509 585
R7666 dvss.n3619 dvss.n510 585
R7667 dvss.n3623 dvss.n510 585
R7668 dvss.n3618 dvss.n3513 585
R7669 dvss.n3513 dvss.n511 585
R7670 dvss.n3563 dvss.n3514 585
R7671 dvss.n3614 dvss.n3517 585
R7672 dvss.n3613 dvss.n3518 585
R7673 dvss.n3567 dvss.n3519 585
R7674 dvss.n3568 dvss.n3526 585
R7675 dvss.n3569 dvss.n3568 585
R7676 dvss.n3606 dvss.n3527 585
R7677 dvss.n3570 dvss.n3527 585
R7678 dvss.n3605 dvss.n3528 585
R7679 dvss.n3573 dvss.n3528 585
R7680 dvss.n3575 dvss.n3529 585
R7681 dvss.n3575 dvss.n3574 585
R7682 dvss.n3576 dvss.n3537 585
R7683 dvss.n3577 dvss.n3576 585
R7684 dvss.n3597 dvss.n3538 585
R7685 dvss.n3580 dvss.n3538 585
R7686 dvss.n3596 dvss.n3539 585
R7687 dvss.n3546 dvss.n3539 585
R7688 dvss.n3545 dvss.n3540 585
R7689 dvss.n3583 dvss.n3545 585
R7690 dvss.n3544 dvss.n376 585
R7691 dvss.n3544 dvss.n3543 585
R7692 dvss.n3891 dvss.n371 585
R7693 dvss.n3895 dvss.n371 585
R7694 dvss.n3890 dvss.n377 585
R7695 dvss.n445 dvss.n377 585
R7696 dvss.n447 dvss.n378 585
R7697 dvss.n447 dvss.n446 585
R7698 dvss.n449 dvss.n448 585
R7699 dvss.n450 dvss.n449 585
R7700 dvss.n443 dvss.n442 585
R7701 dvss.n456 dvss.n443 585
R7702 dvss.n459 dvss.n458 585
R7703 dvss.n458 dvss.n457 585
R7704 dvss.n439 dvss.n389 585
R7705 dvss.n464 dvss.n439 585
R7706 dvss.n3875 dvss.n390 585
R7707 dvss.n3811 dvss.n390 585
R7708 dvss.n3874 dvss.n391 585
R7709 dvss.n3812 dvss.n391 585
R7710 dvss.n430 dvss.n392 585
R7711 dvss.n3870 dvss.n396 585
R7712 dvss.n3869 dvss.n397 585
R7713 dvss.n434 dvss.n398 585
R7714 dvss.n435 dvss.n405 585
R7715 dvss.n3821 dvss.n435 585
R7716 dvss.n3862 dvss.n406 585
R7717 dvss.n3822 dvss.n406 585
R7718 dvss.n3861 dvss.n407 585
R7719 dvss.n3823 dvss.n407 585
R7720 dvss.n425 dvss.n408 585
R7721 dvss.n425 dvss.n424 585
R7722 dvss.n426 dvss.n416 585
R7723 dvss.n3831 dvss.n426 585
R7724 dvss.n3853 dvss.n417 585
R7725 dvss.n3832 dvss.n417 585
R7726 dvss.n3852 dvss.n418 585
R7727 dvss.n3834 dvss.n418 585
R7728 dvss.n3838 dvss.n419 585
R7729 dvss.n3838 dvss.n3837 585
R7730 dvss.n3841 dvss.n3840 585
R7731 dvss.n3840 dvss.n3839 585
R7732 dvss.n347 dvss.n346 585
R7733 dvss.n3932 dvss.n346 585
R7734 dvss.n3939 dvss.n3938 585
R7735 dvss.n3939 dvss.n345 585
R7736 dvss.n3940 dvss.n340 585
R7737 dvss.n3943 dvss.n3940 585
R7738 dvss.n3955 dvss.n341 585
R7739 dvss.n3942 dvss.n341 585
R7740 dvss.n3954 dvss.n330 585
R7741 dvss.n3941 dvss.n330 585
R7742 dvss.n3967 dvss.n331 585
R7743 dvss.n3967 dvss.n3966 585
R7744 dvss.n3968 dvss.n320 585
R7745 dvss.n3969 dvss.n3968 585
R7746 dvss.n3975 dvss.n321 585
R7747 dvss.n3971 dvss.n321 585
R7748 dvss.n3976 dvss.n315 585
R7749 dvss.n316 dvss.n315 585
R7750 dvss.n3982 dvss.n314 585
R7751 dvss.n3982 dvss.n3981 585
R7752 dvss.n3984 dvss.n3983 585
R7753 dvss.n3983 dvss.n306 585
R7754 dvss.n1053 dvss.n1052 585
R7755 dvss.n1050 dvss.n917 585
R7756 dvss.n1049 dvss.n1048 585
R7757 dvss.n1049 dvss.n908 585
R7758 dvss.n1047 dvss.n918 585
R7759 dvss.n1046 dvss.n1045 585
R7760 dvss.n1043 dvss.n922 585
R7761 dvss.n1041 dvss.n1040 585
R7762 dvss.n1039 dvss.n923 585
R7763 dvss.n1038 dvss.n1037 585
R7764 dvss.n1035 dvss.n927 585
R7765 dvss.n1033 dvss.n1032 585
R7766 dvss.n1031 dvss.n928 585
R7767 dvss.n928 dvss.n908 585
R7768 dvss.n966 dvss.n960 585
R7769 dvss.n969 dvss.n968 585
R7770 dvss.n973 dvss.n958 585
R7771 dvss.n958 dvss.n907 585
R7772 dvss.n976 dvss.n975 585
R7773 dvss.n978 dvss.n957 585
R7774 dvss.n981 dvss.n980 585
R7775 dvss.n988 dvss.n955 585
R7776 dvss.n991 dvss.n990 585
R7777 dvss.n993 dvss.n954 585
R7778 dvss.n996 dvss.n995 585
R7779 dvss.n1010 dvss.n952 585
R7780 dvss.n1013 dvss.n1012 585
R7781 dvss.n1013 dvss.n907 585
R7782 dvss.n1230 dvss.n1229 585
R7783 dvss.n1231 dvss.n1230 585
R7784 dvss.n1228 dvss.n1058 585
R7785 dvss.n1058 dvss.n1057 585
R7786 dvss.n1227 dvss.n1226 585
R7787 dvss.n1226 dvss.n1225 585
R7788 dvss.n1062 dvss.n1061 585
R7789 dvss.n1224 dvss.n1062 585
R7790 dvss.n1222 dvss.n1221 585
R7791 dvss.n1223 dvss.n1222 585
R7792 dvss.n1220 dvss.n1064 585
R7793 dvss.n1064 dvss.n1063 585
R7794 dvss.n1219 dvss.n1218 585
R7795 dvss.n1218 dvss.n1217 585
R7796 dvss.n1070 dvss.n1069 585
R7797 dvss.n1216 dvss.n1070 585
R7798 dvss.n1213 dvss.n1212 585
R7799 dvss.n1214 dvss.n1213 585
R7800 dvss.n1211 dvss.n1072 585
R7801 dvss.n1082 dvss.n1072 585
R7802 dvss.n1210 dvss.n1209 585
R7803 dvss.n1209 dvss.n1208 585
R7804 dvss.n1081 dvss.n1080 585
R7805 dvss.n1207 dvss.n1081 585
R7806 dvss.n1205 dvss.n1204 585
R7807 dvss.n1206 dvss.n1205 585
R7808 dvss.n1203 dvss.n1083 585
R7809 dvss.n1095 dvss.n1083 585
R7810 dvss.n1202 dvss.n1201 585
R7811 dvss.n1201 dvss.n1200 585
R7812 dvss.n1094 dvss.n1093 585
R7813 dvss.n1199 dvss.n1094 585
R7814 dvss.n1197 dvss.n1196 585
R7815 dvss.n1198 dvss.n1197 585
R7816 dvss.n1195 dvss.n1097 585
R7817 dvss.n1097 dvss.n1096 585
R7818 dvss.n1194 dvss.n1193 585
R7819 dvss.n1193 dvss.n1192 585
R7820 dvss.n1054 dvss.n913 585
R7821 dvss.n965 dvss.n962 585
R7822 dvss.n2888 dvss.n2887 585
R7823 dvss.n2889 dvss.n2888 585
R7824 dvss.n2392 dvss.n2391 585
R7825 dvss.n2884 dvss.n2393 585
R7826 dvss.n2883 dvss.n2394 585
R7827 dvss.n2396 dvss.n2395 585
R7828 dvss.n2879 dvss.n2397 585
R7829 dvss.n2878 dvss.n2398 585
R7830 dvss.n2400 dvss.n2399 585
R7831 dvss.n2874 dvss.n2401 585
R7832 dvss.n2873 dvss.n2402 585
R7833 dvss.n2407 dvss.n2403 585
R7834 dvss.n2866 dvss.n2408 585
R7835 dvss.n2865 dvss.n2409 585
R7836 dvss.n2411 dvss.n2410 585
R7837 dvss.n2417 dvss.n2416 585
R7838 dvss.n2858 dvss.n2418 585
R7839 dvss.n2857 dvss.n2419 585
R7840 dvss.n2854 dvss.n2420 585
R7841 dvss.n2853 dvss.n2421 585
R7842 dvss.n2423 dvss.n2422 585
R7843 dvss.n2847 dvss.n2427 585
R7844 dvss.n2846 dvss.n2428 585
R7845 dvss.n2430 dvss.n2429 585
R7846 dvss.n2842 dvss.n2431 585
R7847 dvss.n2841 dvss.n2432 585
R7848 dvss.n2434 dvss.n2433 585
R7849 dvss.n2837 dvss.n2435 585
R7850 dvss.n2836 dvss.n2436 585
R7851 dvss.n2440 dvss.n2437 585
R7852 dvss.n2829 dvss.n2441 585
R7853 dvss.n2828 dvss.n2442 585
R7854 dvss.n2444 dvss.n2443 585
R7855 dvss.n2821 dvss.n2446 585
R7856 dvss.n2820 dvss.n2447 585
R7857 dvss.n2449 dvss.n2448 585
R7858 dvss.n2813 dvss.n2450 585
R7859 dvss.n2812 dvss.n2451 585
R7860 dvss.n2453 dvss.n2452 585
R7861 dvss.n2808 dvss.n2454 585
R7862 dvss.n2807 dvss.n2455 585
R7863 dvss.n2460 dvss.n2456 585
R7864 dvss.n2462 dvss.n2461 585
R7865 dvss.n2800 dvss.n2463 585
R7866 dvss.n2799 dvss.n2464 585
R7867 dvss.n2466 dvss.n2465 585
R7868 dvss.n2795 dvss.n2467 585
R7869 dvss.n2794 dvss.n2468 585
R7870 dvss.n2470 dvss.n2469 585
R7871 dvss.n2790 dvss.n2471 585
R7872 dvss.n2789 dvss.n2472 585
R7873 dvss.n2476 dvss.n2473 585
R7874 dvss.n2782 dvss.n2477 585
R7875 dvss.n2781 dvss.n2478 585
R7876 dvss.n2480 dvss.n2479 585
R7877 dvss.n2774 dvss.n2482 585
R7878 dvss.n2773 dvss.n2483 585
R7879 dvss.n2485 dvss.n2484 585
R7880 dvss.n2766 dvss.n2486 585
R7881 dvss.n2765 dvss.n2487 585
R7882 dvss.n2489 dvss.n2488 585
R7883 dvss.n2761 dvss.n2490 585
R7884 dvss.n2760 dvss.n2491 585
R7885 dvss.n2496 dvss.n2492 585
R7886 dvss.n2498 dvss.n2497 585
R7887 dvss.n2753 dvss.n2499 585
R7888 dvss.n2752 dvss.n2500 585
R7889 dvss.n2502 dvss.n2501 585
R7890 dvss.n2748 dvss.n2503 585
R7891 dvss.n2747 dvss.n2504 585
R7892 dvss.n2506 dvss.n2505 585
R7893 dvss.n2743 dvss.n2507 585
R7894 dvss.n2742 dvss.n2508 585
R7895 dvss.n2512 dvss.n2509 585
R7896 dvss.n2735 dvss.n2513 585
R7897 dvss.n2734 dvss.n2514 585
R7898 dvss.n2516 dvss.n2515 585
R7899 dvss.n2727 dvss.n2518 585
R7900 dvss.n2726 dvss.n2519 585
R7901 dvss.n2521 dvss.n2520 585
R7902 dvss.n2719 dvss.n2522 585
R7903 dvss.n2718 dvss.n2523 585
R7904 dvss.n2525 dvss.n2524 585
R7905 dvss.n2714 dvss.n2526 585
R7906 dvss.n2713 dvss.n2527 585
R7907 dvss.n2532 dvss.n2528 585
R7908 dvss.n2534 dvss.n2533 585
R7909 dvss.n2706 dvss.n2535 585
R7910 dvss.n2705 dvss.n2536 585
R7911 dvss.n2538 dvss.n2537 585
R7912 dvss.n2701 dvss.n2539 585
R7913 dvss.n2700 dvss.n2540 585
R7914 dvss.n2542 dvss.n2541 585
R7915 dvss.n2696 dvss.n2543 585
R7916 dvss.n2695 dvss.n2544 585
R7917 dvss.n2548 dvss.n2545 585
R7918 dvss.n2688 dvss.n2549 585
R7919 dvss.n2687 dvss.n2550 585
R7920 dvss.n2552 dvss.n2551 585
R7921 dvss.n2680 dvss.n2554 585
R7922 dvss.n2679 dvss.n2555 585
R7923 dvss.n2557 dvss.n2556 585
R7924 dvss.n2672 dvss.n2558 585
R7925 dvss.n2671 dvss.n2559 585
R7926 dvss.n2561 dvss.n2560 585
R7927 dvss.n2667 dvss.n2562 585
R7928 dvss.n2666 dvss.n2563 585
R7929 dvss.n2568 dvss.n2564 585
R7930 dvss.n2570 dvss.n2569 585
R7931 dvss.n2659 dvss.n2571 585
R7932 dvss.n2658 dvss.n2572 585
R7933 dvss.n2574 dvss.n2573 585
R7934 dvss.n2654 dvss.n2575 585
R7935 dvss.n2653 dvss.n2576 585
R7936 dvss.n2578 dvss.n2577 585
R7937 dvss.n2649 dvss.n2579 585
R7938 dvss.n2648 dvss.n2580 585
R7939 dvss.n2584 dvss.n2581 585
R7940 dvss.n2641 dvss.n2585 585
R7941 dvss.n2640 dvss.n2586 585
R7942 dvss.n2588 dvss.n2587 585
R7943 dvss.n2633 dvss.n2590 585
R7944 dvss.n2632 dvss.n2591 585
R7945 dvss.n2593 dvss.n2592 585
R7946 dvss.n2625 dvss.n2594 585
R7947 dvss.n2624 dvss.n2595 585
R7948 dvss.n2597 dvss.n2596 585
R7949 dvss.n2620 dvss.n2598 585
R7950 dvss.n2619 dvss.n2599 585
R7951 dvss.n2604 dvss.n2600 585
R7952 dvss.n2606 dvss.n2605 585
R7953 dvss.n2612 dvss.n2607 585
R7954 dvss.n2611 dvss.n2608 585
R7955 dvss.n2324 dvss.n2323 585
R7956 dvss.n2892 dvss.n2891 585
R7957 dvss.n2322 dvss.n2321 585
R7958 dvss.n2898 dvss.n2897 585
R7959 dvss.n2899 dvss.n2898 585
R7960 dvss.n2319 dvss.n2318 585
R7961 dvss.n2900 dvss.n2319 585
R7962 dvss.n2903 dvss.n2902 585
R7963 dvss.n2902 dvss.n2901 585
R7964 dvss.n2317 dvss.n2316 585
R7965 dvss.n2316 dvss.n2315 585
R7966 dvss.n2911 dvss.n2910 585
R7967 dvss.n2911 dvss.n2314 585
R7968 dvss.n2912 dvss.n2312 585
R7969 dvss.n2913 dvss.n2912 585
R7970 dvss.n2921 dvss.n2313 585
R7971 dvss.n2914 dvss.n2313 585
R7972 dvss.n2920 dvss.n2917 585
R7973 dvss.n2917 dvss.n2916 585
R7974 dvss.n2307 dvss.n2306 585
R7975 dvss.n2915 dvss.n2306 585
R7976 dvss.n2932 dvss.n2931 585
R7977 dvss.n2933 dvss.n2932 585
R7978 dvss.n2305 dvss.n2304 585
R7979 dvss.n2935 dvss.n2305 585
R7980 dvss.n2938 dvss.n2937 585
R7981 dvss.n2937 dvss.n2936 585
R7982 dvss.n2303 dvss.n2302 585
R7983 dvss.n2302 dvss.n2301 585
R7984 dvss.n2944 dvss.n2943 585
R7985 dvss.n2945 dvss.n2944 585
R7986 dvss.n2300 dvss.n2299 585
R7987 dvss.n2946 dvss.n2300 585
R7988 dvss.n2950 dvss.n2949 585
R7989 dvss.n2949 dvss.n2948 585
R7990 dvss.n2297 dvss.n2296 585
R7991 dvss.n2947 dvss.n2296 585
R7992 dvss.n2960 dvss.n2959 585
R7993 dvss.n2961 dvss.n2960 585
R7994 dvss.n2295 dvss.n2294 585
R7995 dvss.n2962 dvss.n2295 585
R7996 dvss.n2965 dvss.n2964 585
R7997 dvss.n2964 dvss.n2963 585
R7998 dvss.n2293 dvss.n2292 585
R7999 dvss.n2292 dvss.n2291 585
R8000 dvss.n2971 dvss.n2970 585
R8001 dvss.n2972 dvss.n2971 585
R8002 dvss.n2290 dvss.n2289 585
R8003 dvss.n2973 dvss.n2290 585
R8004 dvss.n2977 dvss.n2976 585
R8005 dvss.n2976 dvss.n2975 585
R8006 dvss.n2212 dvss.n2210 585
R8007 dvss.n2974 dvss.n2210 585
R8008 dvss.n2985 dvss.n2984 585
R8009 dvss.n2986 dvss.n2985 585
R8010 dvss.n2213 dvss.n2211 585
R8011 dvss.n2224 dvss.n2211 585
R8012 dvss.n2227 dvss.n2226 585
R8013 dvss.n2226 dvss.n2225 585
R8014 dvss.n2221 dvss.n2220 585
R8015 dvss.n2220 dvss.n2219 585
R8016 dvss.n2236 dvss.n2235 585
R8017 dvss.n2237 dvss.n2236 585
R8018 dvss.n2222 dvss.n2218 585
R8019 dvss.n2238 dvss.n2218 585
R8020 dvss.n2240 dvss.n2217 585
R8021 dvss.n2240 dvss.n2239 585
R8022 dvss.n2283 dvss.n2241 585
R8023 dvss.n2251 dvss.n2241 585
R8024 dvss.n2282 dvss.n2242 585
R8025 dvss.n2252 dvss.n2242 585
R8026 dvss.n2253 dvss.n2243 585
R8027 dvss.n2254 dvss.n2253 585
R8028 dvss.n2278 dvss.n2244 585
R8029 dvss.n2255 dvss.n2244 585
R8030 dvss.n2277 dvss.n2245 585
R8031 dvss.n2256 dvss.n2245 585
R8032 dvss.n2249 dvss.n2246 585
R8033 dvss.n2257 dvss.n2249 585
R8034 dvss.n2270 dvss.n2269 585
R8035 dvss.n2269 dvss.n2268 585
R8036 dvss.n2250 dvss.n259 585
R8037 dvss.n2267 dvss.n2250 585
R8038 dvss.n4131 dvss.n260 585
R8039 dvss.n2266 dvss.n260 585
R8040 dvss.n4130 dvss.n261 585
R8041 dvss.n2265 dvss.n261 585
R8042 dvss.n2263 dvss.n262 585
R8043 dvss.n2264 dvss.n2263 585
R8044 dvss.n4126 dvss.n263 585
R8045 dvss.n2262 dvss.n263 585
R8046 dvss.n4125 dvss.n264 585
R8047 dvss.n2261 dvss.n264 585
R8048 dvss.n2259 dvss.n265 585
R8049 dvss.n2260 dvss.n2259 585
R8050 dvss.n4121 dvss.n266 585
R8051 dvss.n2258 dvss.n266 585
R8052 dvss.n4120 dvss.n267 585
R8053 dvss.n355 dvss.n267 585
R8054 dvss.n369 dvss.n268 585
R8055 dvss.n370 dvss.n369 585
R8056 dvss.n368 dvss.n367 585
R8057 dvss.n368 dvss.n353 585
R8058 dvss.n357 dvss.n356 585
R8059 dvss.n356 dvss.n354 585
R8060 dvss.n361 dvss.n350 585
R8061 dvss.n3900 dvss.n351 585
R8062 dvss.n3901 dvss.n272 585
R8063 dvss.n3902 dvss.n3901 585
R8064 dvss.n4110 dvss.n273 585
R8065 dvss.n3903 dvss.n273 585
R8066 dvss.n4109 dvss.n274 585
R8067 dvss.n3904 dvss.n274 585
R8068 dvss.n3905 dvss.n275 585
R8069 dvss.n3906 dvss.n3905 585
R8070 dvss.n4105 dvss.n276 585
R8071 dvss.n3907 dvss.n276 585
R8072 dvss.n4104 dvss.n277 585
R8073 dvss.n3908 dvss.n277 585
R8074 dvss.n3910 dvss.n278 585
R8075 dvss.n3910 dvss.n3909 585
R8076 dvss.n3911 dvss.n282 585
R8077 dvss.n3912 dvss.n3911 585
R8078 dvss.n4097 dvss.n283 585
R8079 dvss.n3913 dvss.n283 585
R8080 dvss.n4096 dvss.n284 585
R8081 dvss.n3914 dvss.n284 585
R8082 dvss.n3915 dvss.n285 585
R8083 dvss.n3916 dvss.n3915 585
R8084 dvss.n4092 dvss.n286 585
R8085 dvss.n3917 dvss.n286 585
R8086 dvss.n4091 dvss.n287 585
R8087 dvss.n3918 dvss.n287 585
R8088 dvss.n3919 dvss.n288 585
R8089 dvss.n3920 dvss.n3919 585
R8090 dvss.n4087 dvss.n289 585
R8091 dvss.n3921 dvss.n289 585
R8092 dvss.n4086 dvss.n290 585
R8093 dvss.n3922 dvss.n290 585
R8094 dvss.n3927 dvss.n291 585
R8095 dvss.n3928 dvss.n3927 585
R8096 dvss.n4079 dvss.n294 585
R8097 dvss.n3930 dvss.n294 585
R8098 dvss.n4078 dvss.n295 585
R8099 dvss.n3929 dvss.n295 585
R8100 dvss.n3923 dvss.n296 585
R8101 dvss.n4071 dvss.n298 585
R8102 dvss.n4070 dvss.n299 585
R8103 dvss.n327 dvss.n300 585
R8104 dvss.n328 dvss.n327 585
R8105 dvss.n4063 dvss.n301 585
R8106 dvss.n326 dvss.n301 585
R8107 dvss.n4062 dvss.n302 585
R8108 dvss.n325 dvss.n302 585
R8109 dvss.n304 dvss.n303 585
R8110 dvss.n305 dvss.n304 585
R8111 dvss.n4058 dvss.n4057 585
R8112 dvss.n4057 dvss.n4056 585
R8113 dvss.n4055 dvss.n306 583.256
R8114 dvss.n133 dvss.t713 575.611
R8115 dvss.t416 dvss.n174 568.053
R8116 dvss.n432 dvss.n429 564.282
R8117 dvss.n3565 dvss.n3562 564.282
R8118 dvss.n3419 dvss.n563 564.282
R8119 dvss.n3294 dvss.n3292 564.282
R8120 dvss.n3166 dvss.n687 564.282
R8121 dvss.n1865 dvss.n1862 564.282
R8122 dvss.n1688 dvss.n796 564.282
R8123 dvss.n1390 dvss.n1387 564.282
R8124 dvss.n1233 dvss.n912 561.928
R8125 dvss.n1233 dvss.n1232 561.928
R8126 dvss.n1230 dvss.n1058 539.294
R8127 dvss.n1226 dvss.n1058 539.294
R8128 dvss.n1226 dvss.n1062 539.294
R8129 dvss.n1222 dvss.n1062 539.294
R8130 dvss.n1222 dvss.n1064 539.294
R8131 dvss.n1218 dvss.n1064 539.294
R8132 dvss.n1218 dvss.n1070 539.294
R8133 dvss.n1213 dvss.n1070 539.294
R8134 dvss.n1213 dvss.n1072 539.294
R8135 dvss.n1209 dvss.n1072 539.294
R8136 dvss.n1209 dvss.n1081 539.294
R8137 dvss.n1205 dvss.n1081 539.294
R8138 dvss.n1205 dvss.n1083 539.294
R8139 dvss.n1201 dvss.n1083 539.294
R8140 dvss.n1201 dvss.n1094 539.294
R8141 dvss.n1197 dvss.n1094 539.294
R8142 dvss.n1193 dvss.n1097 539.294
R8143 dvss.n1193 dvss.n1107 539.294
R8144 dvss.n1189 dvss.n1107 539.294
R8145 dvss.n1189 dvss.n1108 539.294
R8146 dvss.n1185 dvss.n1108 539.294
R8147 dvss.n1185 dvss.n1114 539.294
R8148 dvss.n1181 dvss.n1114 539.294
R8149 dvss.n1181 dvss.n1116 539.294
R8150 dvss.n1177 dvss.n1116 539.294
R8151 dvss.n1177 dvss.n1121 539.294
R8152 dvss.n1173 dvss.n1121 539.294
R8153 dvss.n1173 dvss.n1126 539.294
R8154 dvss.n1169 dvss.n1126 539.294
R8155 dvss.n1169 dvss.n1149 539.294
R8156 dvss.n1165 dvss.n1149 539.294
R8157 dvss.n1165 dvss.n1151 539.294
R8158 dvss.n1151 dvss.n851 539.294
R8159 dvss.n1495 dvss.n851 539.294
R8160 dvss.n1495 dvss.n848 539.294
R8161 dvss.n1502 dvss.n848 539.294
R8162 dvss.n1506 dvss.n847 539.294
R8163 dvss.n1514 dvss.n844 539.294
R8164 dvss.n1514 dvss.n842 539.294
R8165 dvss.n1518 dvss.n842 539.294
R8166 dvss.n1518 dvss.n836 539.294
R8167 dvss.n1529 dvss.n836 539.294
R8168 dvss.n1529 dvss.n834 539.294
R8169 dvss.n1534 dvss.n834 539.294
R8170 dvss.n1534 dvss.n826 539.294
R8171 dvss.n1544 dvss.n826 539.294
R8172 dvss.n1544 dvss.n825 539.294
R8173 dvss.n1549 dvss.n825 539.294
R8174 dvss.n1549 dvss.n818 539.294
R8175 dvss.n1559 dvss.n818 539.294
R8176 dvss.n1559 dvss.n817 539.294
R8177 dvss.n1563 dvss.n817 539.294
R8178 dvss.n1563 dvss.n812 539.294
R8179 dvss.n1672 dvss.n812 539.294
R8180 dvss.n1672 dvss.n813 539.294
R8181 dvss.n1567 dvss.n813 539.294
R8182 dvss.n1595 dvss.n1568 539.294
R8183 dvss.n1571 dvss.n1570 539.294
R8184 dvss.n1602 dvss.n1571 539.294
R8185 dvss.n1603 dvss.n1602 539.294
R8186 dvss.n1603 dvss.n1576 539.294
R8187 dvss.n1577 dvss.n1576 539.294
R8188 dvss.n1594 dvss.n1577 539.294
R8189 dvss.n1594 dvss.n1582 539.294
R8190 dvss.n1583 dvss.n1582 539.294
R8191 dvss.n1612 dvss.n1583 539.294
R8192 dvss.n1612 dvss.n1586 539.294
R8193 dvss.n1587 dvss.n1586 539.294
R8194 dvss.n1617 dvss.n1587 539.294
R8195 dvss.n1618 dvss.n1617 539.294
R8196 dvss.n1618 dvss.n1593 539.294
R8197 dvss.n1622 dvss.n1593 539.294
R8198 dvss.n1622 dvss.n742 539.294
R8199 dvss.n1970 dvss.n742 539.294
R8200 dvss.n1970 dvss.n739 539.294
R8201 dvss.n1977 dvss.n739 539.294
R8202 dvss.n1981 dvss.n738 539.294
R8203 dvss.n1989 dvss.n735 539.294
R8204 dvss.n1989 dvss.n733 539.294
R8205 dvss.n1993 dvss.n733 539.294
R8206 dvss.n1993 dvss.n727 539.294
R8207 dvss.n2004 dvss.n727 539.294
R8208 dvss.n2004 dvss.n725 539.294
R8209 dvss.n2009 dvss.n725 539.294
R8210 dvss.n2009 dvss.n717 539.294
R8211 dvss.n2019 dvss.n717 539.294
R8212 dvss.n2019 dvss.n716 539.294
R8213 dvss.n2024 dvss.n716 539.294
R8214 dvss.n2024 dvss.n709 539.294
R8215 dvss.n2034 dvss.n709 539.294
R8216 dvss.n2034 dvss.n708 539.294
R8217 dvss.n2038 dvss.n708 539.294
R8218 dvss.n2038 dvss.n703 539.294
R8219 dvss.n3150 dvss.n703 539.294
R8220 dvss.n3150 dvss.n704 539.294
R8221 dvss.n2042 dvss.n704 539.294
R8222 dvss.n2144 dvss.n2043 539.294
R8223 dvss.n2046 dvss.n2045 539.294
R8224 dvss.n2151 dvss.n2046 539.294
R8225 dvss.n2152 dvss.n2151 539.294
R8226 dvss.n2152 dvss.n2051 539.294
R8227 dvss.n2052 dvss.n2051 539.294
R8228 dvss.n2143 dvss.n2052 539.294
R8229 dvss.n2143 dvss.n2057 539.294
R8230 dvss.n2058 dvss.n2057 539.294
R8231 dvss.n2161 dvss.n2058 539.294
R8232 dvss.n2161 dvss.n2061 539.294
R8233 dvss.n2062 dvss.n2061 539.294
R8234 dvss.n2166 dvss.n2062 539.294
R8235 dvss.n2167 dvss.n2166 539.294
R8236 dvss.n2167 dvss.n2068 539.294
R8237 dvss.n2069 dvss.n2068 539.294
R8238 dvss.n2171 dvss.n2069 539.294
R8239 dvss.n2171 dvss.n2071 539.294
R8240 dvss.n2072 dvss.n2071 539.294
R8241 dvss.n2140 dvss.n2072 539.294
R8242 dvss.n2075 dvss.n2074 539.294
R8243 dvss.n2138 dvss.n2077 539.294
R8244 dvss.n2078 dvss.n2077 539.294
R8245 dvss.n2179 dvss.n2078 539.294
R8246 dvss.n2179 dvss.n2082 539.294
R8247 dvss.n2083 dvss.n2082 539.294
R8248 dvss.n2137 dvss.n2083 539.294
R8249 dvss.n2137 dvss.n2088 539.294
R8250 dvss.n2089 dvss.n2088 539.294
R8251 dvss.n2186 dvss.n2089 539.294
R8252 dvss.n2186 dvss.n2092 539.294
R8253 dvss.n2093 dvss.n2092 539.294
R8254 dvss.n2191 dvss.n2093 539.294
R8255 dvss.n2192 dvss.n2191 539.294
R8256 dvss.n2192 dvss.n2099 539.294
R8257 dvss.n2100 dvss.n2099 539.294
R8258 dvss.n2196 dvss.n2100 539.294
R8259 dvss.n2196 dvss.n2102 539.294
R8260 dvss.n2103 dvss.n2102 539.294
R8261 dvss.n2134 dvss.n2103 539.294
R8262 dvss.n2106 dvss.n2105 539.294
R8263 dvss.n2132 dvss.n2108 539.294
R8264 dvss.n2109 dvss.n2108 539.294
R8265 dvss.n2204 dvss.n2109 539.294
R8266 dvss.n2204 dvss.n2113 539.294
R8267 dvss.n2114 dvss.n2113 539.294
R8268 dvss.n2131 dvss.n2114 539.294
R8269 dvss.n2131 dvss.n2119 539.294
R8270 dvss.n2120 dvss.n2119 539.294
R8271 dvss.n2990 dvss.n2120 539.294
R8272 dvss.n2990 dvss.n2123 539.294
R8273 dvss.n2124 dvss.n2123 539.294
R8274 dvss.n2995 dvss.n2124 539.294
R8275 dvss.n2996 dvss.n2995 539.294
R8276 dvss.n2996 dvss.n2130 539.294
R8277 dvss.n3000 dvss.n2130 539.294
R8278 dvss.n3000 dvss.n506 539.294
R8279 dvss.n3628 dvss.n506 539.294
R8280 dvss.n3628 dvss.n503 539.294
R8281 dvss.n3635 dvss.n503 539.294
R8282 dvss.n3639 dvss.n502 539.294
R8283 dvss.n3647 dvss.n499 539.294
R8284 dvss.n3647 dvss.n497 539.294
R8285 dvss.n3651 dvss.n497 539.294
R8286 dvss.n3651 dvss.n491 539.294
R8287 dvss.n3662 dvss.n491 539.294
R8288 dvss.n3662 dvss.n489 539.294
R8289 dvss.n3667 dvss.n489 539.294
R8290 dvss.n3667 dvss.n481 539.294
R8291 dvss.n3677 dvss.n481 539.294
R8292 dvss.n3677 dvss.n480 539.294
R8293 dvss.n3682 dvss.n480 539.294
R8294 dvss.n3682 dvss.n473 539.294
R8295 dvss.n3692 dvss.n473 539.294
R8296 dvss.n3692 dvss.n472 539.294
R8297 dvss.n3696 dvss.n472 539.294
R8298 dvss.n3696 dvss.n467 539.294
R8299 dvss.n3807 dvss.n467 539.294
R8300 dvss.n3807 dvss.n468 539.294
R8301 dvss.n3700 dvss.n468 539.294
R8302 dvss.n3717 dvss.n3701 539.294
R8303 dvss.n3704 dvss.n3703 539.294
R8304 dvss.n3724 dvss.n3704 539.294
R8305 dvss.n3725 dvss.n3724 539.294
R8306 dvss.n3725 dvss.n3709 539.294
R8307 dvss.n3710 dvss.n3709 539.294
R8308 dvss.n3716 dvss.n3710 539.294
R8309 dvss.n3716 dvss.n3715 539.294
R8310 dvss.n3732 dvss.n3715 539.294
R8311 dvss.n3744 dvss.n3732 539.294
R8312 dvss.n3744 dvss.n3735 539.294
R8313 dvss.n3736 dvss.n3735 539.294
R8314 dvss.n3749 dvss.n3736 539.294
R8315 dvss.n3750 dvss.n3749 539.294
R8316 dvss.n3750 dvss.n3742 539.294
R8317 dvss.n3743 dvss.n3742 539.294
R8318 dvss.n3755 dvss.n3743 539.294
R8319 dvss.n3755 dvss.n309 539.294
R8320 dvss.n4052 dvss.n309 539.294
R8321 dvss.n4052 dvss.n310 539.294
R8322 dvss.n966 dvss.n965 539.294
R8323 dvss.n968 dvss.n958 539.294
R8324 dvss.n976 dvss.n958 539.294
R8325 dvss.n980 dvss.n978 539.294
R8326 dvss.n991 dvss.n955 539.294
R8327 dvss.n995 dvss.n993 539.294
R8328 dvss.n1013 dvss.n952 539.294
R8329 dvss.n1014 dvss.n1013 539.294
R8330 dvss.n1016 dvss.n951 539.294
R8331 dvss.n951 dvss.n950 539.294
R8332 dvss.n937 dvss.n899 539.294
R8333 dvss.n1246 dvss.n899 539.294
R8334 dvss.n1246 dvss.n895 539.294
R8335 dvss.n1259 dvss.n895 539.294
R8336 dvss.n1260 dvss.n1259 539.294
R8337 dvss.n1260 dvss.n889 539.294
R8338 dvss.n889 dvss.n884 539.294
R8339 dvss.n1283 dvss.n884 539.294
R8340 dvss.n1284 dvss.n1283 539.294
R8341 dvss.n1284 dvss.n880 539.294
R8342 dvss.n880 dvss.n874 539.294
R8343 dvss.n1308 dvss.n874 539.294
R8344 dvss.n1309 dvss.n1308 539.294
R8345 dvss.n1309 dvss.n873 539.294
R8346 dvss.n1314 dvss.n873 539.294
R8347 dvss.n1314 dvss.n856 539.294
R8348 dvss.n1489 dvss.n856 539.294
R8349 dvss.n1489 dvss.n857 539.294
R8350 dvss.n1396 dvss.n857 539.294
R8351 dvss.n1395 dvss.n1394 539.294
R8352 dvss.n1402 dvss.n1400 539.294
R8353 dvss.n1402 dvss.n1385 539.294
R8354 dvss.n1406 dvss.n1385 539.294
R8355 dvss.n1407 dvss.n1406 539.294
R8356 dvss.n1412 dvss.n1407 539.294
R8357 dvss.n1412 dvss.n1381 539.294
R8358 dvss.n1417 dvss.n1381 539.294
R8359 dvss.n1418 dvss.n1417 539.294
R8360 dvss.n1418 dvss.n1379 539.294
R8361 dvss.n1425 dvss.n1379 539.294
R8362 dvss.n1426 dvss.n1425 539.294
R8363 dvss.n1426 dvss.n1376 539.294
R8364 dvss.n1432 dvss.n1376 539.294
R8365 dvss.n1433 dvss.n1432 539.294
R8366 dvss.n1433 dvss.n808 539.294
R8367 dvss.n1677 dvss.n808 539.294
R8368 dvss.n1677 dvss.n800 539.294
R8369 dvss.n1706 dvss.n800 539.294
R8370 dvss.n1706 dvss.n801 539.294
R8371 dvss.n1697 dvss.n1694 539.294
R8372 dvss.n1695 dvss.n790 539.294
R8373 dvss.n1721 dvss.n790 539.294
R8374 dvss.n1721 dvss.n786 539.294
R8375 dvss.n1734 dvss.n786 539.294
R8376 dvss.n1735 dvss.n1734 539.294
R8377 dvss.n1735 dvss.n780 539.294
R8378 dvss.n780 dvss.n775 539.294
R8379 dvss.n1758 dvss.n775 539.294
R8380 dvss.n1759 dvss.n1758 539.294
R8381 dvss.n1759 dvss.n771 539.294
R8382 dvss.n771 dvss.n765 539.294
R8383 dvss.n1783 dvss.n765 539.294
R8384 dvss.n1784 dvss.n1783 539.294
R8385 dvss.n1784 dvss.n764 539.294
R8386 dvss.n1789 dvss.n764 539.294
R8387 dvss.n1789 dvss.n747 539.294
R8388 dvss.n1964 dvss.n747 539.294
R8389 dvss.n1964 dvss.n748 539.294
R8390 dvss.n1871 dvss.n748 539.294
R8391 dvss.n1870 dvss.n1869 539.294
R8392 dvss.n1877 dvss.n1875 539.294
R8393 dvss.n1877 dvss.n1860 539.294
R8394 dvss.n1881 dvss.n1860 539.294
R8395 dvss.n1882 dvss.n1881 539.294
R8396 dvss.n1887 dvss.n1882 539.294
R8397 dvss.n1887 dvss.n1856 539.294
R8398 dvss.n1892 dvss.n1856 539.294
R8399 dvss.n1893 dvss.n1892 539.294
R8400 dvss.n1893 dvss.n1854 539.294
R8401 dvss.n1900 dvss.n1854 539.294
R8402 dvss.n1901 dvss.n1900 539.294
R8403 dvss.n1901 dvss.n1851 539.294
R8404 dvss.n1907 dvss.n1851 539.294
R8405 dvss.n1908 dvss.n1907 539.294
R8406 dvss.n1908 dvss.n699 539.294
R8407 dvss.n3155 dvss.n699 539.294
R8408 dvss.n3155 dvss.n691 539.294
R8409 dvss.n3184 dvss.n691 539.294
R8410 dvss.n3184 dvss.n692 539.294
R8411 dvss.n3175 dvss.n3172 539.294
R8412 dvss.n3173 dvss.n681 539.294
R8413 dvss.n3199 dvss.n681 539.294
R8414 dvss.n3199 dvss.n677 539.294
R8415 dvss.n3212 dvss.n677 539.294
R8416 dvss.n3213 dvss.n3212 539.294
R8417 dvss.n3213 dvss.n671 539.294
R8418 dvss.n671 dvss.n666 539.294
R8419 dvss.n3236 dvss.n666 539.294
R8420 dvss.n3237 dvss.n3236 539.294
R8421 dvss.n3237 dvss.n662 539.294
R8422 dvss.n662 dvss.n656 539.294
R8423 dvss.n3261 dvss.n656 539.294
R8424 dvss.n3262 dvss.n3261 539.294
R8425 dvss.n3262 dvss.n655 539.294
R8426 dvss.n3268 dvss.n655 539.294
R8427 dvss.n3268 dvss.n639 539.294
R8428 dvss.n3285 dvss.n639 539.294
R8429 dvss.n3285 dvss.n633 539.294
R8430 dvss.n3304 dvss.n633 539.294
R8431 dvss.n632 dvss.n629 539.294
R8432 dvss.n3308 dvss.n622 539.294
R8433 dvss.n3321 dvss.n622 539.294
R8434 dvss.n3321 dvss.n619 539.294
R8435 dvss.n3328 dvss.n619 539.294
R8436 dvss.n3328 dvss.n612 539.294
R8437 dvss.n3347 dvss.n612 539.294
R8438 dvss.n3347 dvss.n607 539.294
R8439 dvss.n3352 dvss.n607 539.294
R8440 dvss.n3352 dvss.n601 539.294
R8441 dvss.n3364 dvss.n601 539.294
R8442 dvss.n3364 dvss.n596 539.294
R8443 dvss.n3378 dvss.n596 539.294
R8444 dvss.n3378 dvss.n592 539.294
R8445 dvss.n3385 dvss.n592 539.294
R8446 dvss.n3385 dvss.n593 539.294
R8447 dvss.n593 dvss.n581 539.294
R8448 dvss.n581 dvss.n574 539.294
R8449 dvss.n3406 dvss.n574 539.294
R8450 dvss.n3407 dvss.n3406 539.294
R8451 dvss.n3411 dvss.n570 539.294
R8452 dvss.n571 dvss.n560 539.294
R8453 dvss.n560 dvss.n555 539.294
R8454 dvss.n3443 dvss.n555 539.294
R8455 dvss.n3444 dvss.n3443 539.294
R8456 dvss.n3444 dvss.n544 539.294
R8457 dvss.n3463 dvss.n544 539.294
R8458 dvss.n3463 dvss.n540 539.294
R8459 dvss.n3468 dvss.n540 539.294
R8460 dvss.n3469 dvss.n3468 539.294
R8461 dvss.n3469 dvss.n536 539.294
R8462 dvss.n536 dvss.n530 539.294
R8463 dvss.n3493 dvss.n530 539.294
R8464 dvss.n3494 dvss.n3493 539.294
R8465 dvss.n3494 dvss.n529 539.294
R8466 dvss.n3499 dvss.n529 539.294
R8467 dvss.n3499 dvss.n512 539.294
R8468 dvss.n3622 dvss.n512 539.294
R8469 dvss.n3622 dvss.n513 539.294
R8470 dvss.n3558 dvss.n513 539.294
R8471 dvss.n3557 dvss.n3556 539.294
R8472 dvss.n3554 dvss.n3553 539.294
R8473 dvss.n3571 dvss.n3553 539.294
R8474 dvss.n3572 dvss.n3571 539.294
R8475 dvss.n3572 dvss.n3547 539.294
R8476 dvss.n3578 dvss.n3547 539.294
R8477 dvss.n3579 dvss.n3578 539.294
R8478 dvss.n3579 dvss.n3542 539.294
R8479 dvss.n3584 dvss.n3542 539.294
R8480 dvss.n3584 dvss.n372 539.294
R8481 dvss.n3894 dvss.n372 539.294
R8482 dvss.n3894 dvss.n373 539.294
R8483 dvss.n444 dvss.n373 539.294
R8484 dvss.n451 dvss.n444 539.294
R8485 dvss.n455 dvss.n451 539.294
R8486 dvss.n455 dvss.n440 539.294
R8487 dvss.n463 dvss.n440 539.294
R8488 dvss.n463 dvss.n438 539.294
R8489 dvss.n3813 dvss.n438 539.294
R8490 dvss.n3814 dvss.n3813 539.294
R8491 dvss.n437 dvss.n436 539.294
R8492 dvss.n3820 dvss.n3818 539.294
R8493 dvss.n3820 dvss.n427 539.294
R8494 dvss.n3824 dvss.n427 539.294
R8495 dvss.n3825 dvss.n3824 539.294
R8496 dvss.n3830 dvss.n3825 539.294
R8497 dvss.n3830 dvss.n423 539.294
R8498 dvss.n3835 dvss.n423 539.294
R8499 dvss.n3836 dvss.n3835 539.294
R8500 dvss.n3836 dvss.n349 539.294
R8501 dvss.n3933 dvss.n349 539.294
R8502 dvss.n3933 dvss.n343 539.294
R8503 dvss.n3944 dvss.n343 539.294
R8504 dvss.n3944 dvss.n344 539.294
R8505 dvss.n344 dvss.n332 539.294
R8506 dvss.n3965 dvss.n332 539.294
R8507 dvss.n3965 dvss.n324 539.294
R8508 dvss.n3972 dvss.n324 539.294
R8509 dvss.n3972 dvss.n317 539.294
R8510 dvss.n3980 dvss.n317 539.294
R8511 dvss.n3980 dvss.n318 539.294
R8512 dvss.n1052 dvss.n913 539.294
R8513 dvss.n1050 dvss.n1049 539.294
R8514 dvss.n1049 dvss.n918 539.294
R8515 dvss.n1045 dvss.n1043 539.294
R8516 dvss.n1041 dvss.n923 539.294
R8517 dvss.n1037 dvss.n1035 539.294
R8518 dvss.n1033 dvss.n928 539.294
R8519 dvss.n931 dvss.n928 539.294
R8520 dvss.n941 dvss.n931 539.294
R8521 dvss.n1235 dvss.n904 539.294
R8522 dvss.n1235 dvss.n898 539.294
R8523 dvss.n1249 dvss.n898 539.294
R8524 dvss.n1249 dvss.n892 539.294
R8525 dvss.n1262 dvss.n892 539.294
R8526 dvss.n1262 dvss.n886 539.294
R8527 dvss.n1278 dvss.n886 539.294
R8528 dvss.n1278 dvss.n883 539.294
R8529 dvss.n1286 dvss.n883 539.294
R8530 dvss.n1286 dvss.n877 539.294
R8531 dvss.n1305 dvss.n877 539.294
R8532 dvss.n1306 dvss.n1305 539.294
R8533 dvss.n1306 dvss.n870 539.294
R8534 dvss.n871 dvss.n870 539.294
R8535 dvss.n1312 dvss.n871 539.294
R8536 dvss.n1312 dvss.n862 539.294
R8537 dvss.n862 dvss.n854 539.294
R8538 dvss.n1328 dvss.n854 539.294
R8539 dvss.n1388 dvss.n1328 539.294
R8540 dvss.n1333 dvss.n1332 539.294
R8541 dvss.n1393 dvss.n1392 539.294
R8542 dvss.n1393 dvss.n1342 539.294
R8543 dvss.n1343 dvss.n1342 539.294
R8544 dvss.n1383 dvss.n1343 539.294
R8545 dvss.n1384 dvss.n1383 539.294
R8546 dvss.n1384 dvss.n1353 539.294
R8547 dvss.n1354 dvss.n1353 539.294
R8548 dvss.n1420 dvss.n1354 539.294
R8549 dvss.n1421 dvss.n1420 539.294
R8550 dvss.n1421 dvss.n1362 539.294
R8551 dvss.n1363 dvss.n1362 539.294
R8552 dvss.n1429 dvss.n1363 539.294
R8553 dvss.n1430 dvss.n1429 539.294
R8554 dvss.n1430 dvss.n1375 539.294
R8555 dvss.n1436 dvss.n1375 539.294
R8556 dvss.n1436 dvss.n809 539.294
R8557 dvss.n809 dvss.n805 539.294
R8558 dvss.n805 dvss.n799 539.294
R8559 dvss.n1685 dvss.n799 539.294
R8560 dvss.n1690 dvss.n1686 539.294
R8561 dvss.n1710 dvss.n795 539.294
R8562 dvss.n1710 dvss.n789 539.294
R8563 dvss.n1724 dvss.n789 539.294
R8564 dvss.n1724 dvss.n783 539.294
R8565 dvss.n1737 dvss.n783 539.294
R8566 dvss.n1737 dvss.n777 539.294
R8567 dvss.n1753 dvss.n777 539.294
R8568 dvss.n1753 dvss.n774 539.294
R8569 dvss.n1761 dvss.n774 539.294
R8570 dvss.n1761 dvss.n768 539.294
R8571 dvss.n1780 dvss.n768 539.294
R8572 dvss.n1781 dvss.n1780 539.294
R8573 dvss.n1781 dvss.n761 539.294
R8574 dvss.n762 dvss.n761 539.294
R8575 dvss.n1787 dvss.n762 539.294
R8576 dvss.n1787 dvss.n753 539.294
R8577 dvss.n753 dvss.n745 539.294
R8578 dvss.n1803 dvss.n745 539.294
R8579 dvss.n1863 dvss.n1803 539.294
R8580 dvss.n1808 dvss.n1807 539.294
R8581 dvss.n1868 dvss.n1867 539.294
R8582 dvss.n1868 dvss.n1817 539.294
R8583 dvss.n1818 dvss.n1817 539.294
R8584 dvss.n1858 dvss.n1818 539.294
R8585 dvss.n1859 dvss.n1858 539.294
R8586 dvss.n1859 dvss.n1828 539.294
R8587 dvss.n1829 dvss.n1828 539.294
R8588 dvss.n1895 dvss.n1829 539.294
R8589 dvss.n1896 dvss.n1895 539.294
R8590 dvss.n1896 dvss.n1837 539.294
R8591 dvss.n1838 dvss.n1837 539.294
R8592 dvss.n1904 dvss.n1838 539.294
R8593 dvss.n1905 dvss.n1904 539.294
R8594 dvss.n1905 dvss.n1850 539.294
R8595 dvss.n1911 dvss.n1850 539.294
R8596 dvss.n1911 dvss.n700 539.294
R8597 dvss.n700 dvss.n696 539.294
R8598 dvss.n696 dvss.n690 539.294
R8599 dvss.n3163 dvss.n690 539.294
R8600 dvss.n3168 dvss.n3164 539.294
R8601 dvss.n3188 dvss.n686 539.294
R8602 dvss.n3188 dvss.n680 539.294
R8603 dvss.n3202 dvss.n680 539.294
R8604 dvss.n3202 dvss.n674 539.294
R8605 dvss.n3215 dvss.n674 539.294
R8606 dvss.n3215 dvss.n668 539.294
R8607 dvss.n3231 dvss.n668 539.294
R8608 dvss.n3231 dvss.n665 539.294
R8609 dvss.n3239 dvss.n665 539.294
R8610 dvss.n3239 dvss.n659 539.294
R8611 dvss.n3258 dvss.n659 539.294
R8612 dvss.n3259 dvss.n3258 539.294
R8613 dvss.n3259 dvss.n652 539.294
R8614 dvss.n653 dvss.n652 539.294
R8615 dvss.n3265 dvss.n653 539.294
R8616 dvss.n3265 dvss.n644 539.294
R8617 dvss.n644 dvss.n637 539.294
R8618 dvss.n3288 dvss.n637 539.294
R8619 dvss.n3289 dvss.n3288 539.294
R8620 dvss.n3296 dvss.n3290 539.294
R8621 dvss.n3291 dvss.n627 539.294
R8622 dvss.n627 dvss.n620 539.294
R8623 dvss.n3324 dvss.n620 539.294
R8624 dvss.n3325 dvss.n3324 539.294
R8625 dvss.n3325 dvss.n615 539.294
R8626 dvss.n615 dvss.n611 539.294
R8627 dvss.n611 dvss.n610 539.294
R8628 dvss.n610 dvss.n605 539.294
R8629 dvss.n605 dvss.n599 539.294
R8630 dvss.n3366 dvss.n599 539.294
R8631 dvss.n3367 dvss.n3366 539.294
R8632 dvss.n3367 dvss.n595 539.294
R8633 dvss.n595 dvss.n589 539.294
R8634 dvss.n590 dvss.n589 539.294
R8635 dvss.n3381 dvss.n590 539.294
R8636 dvss.n3381 dvss.n577 539.294
R8637 dvss.n3403 dvss.n577 539.294
R8638 dvss.n3403 dvss.n565 539.294
R8639 dvss.n3417 dvss.n565 539.294
R8640 dvss.n564 dvss.n562 539.294
R8641 dvss.n3421 dvss.n557 539.294
R8642 dvss.n3440 dvss.n557 539.294
R8643 dvss.n3440 dvss.n552 539.294
R8644 dvss.n3446 dvss.n552 539.294
R8645 dvss.n3446 dvss.n553 539.294
R8646 dvss.n553 dvss.n543 539.294
R8647 dvss.n548 dvss.n543 539.294
R8648 dvss.n548 dvss.n539 539.294
R8649 dvss.n3471 dvss.n539 539.294
R8650 dvss.n3471 dvss.n533 539.294
R8651 dvss.n3490 dvss.n533 539.294
R8652 dvss.n3491 dvss.n3490 539.294
R8653 dvss.n3491 dvss.n526 539.294
R8654 dvss.n527 dvss.n526 539.294
R8655 dvss.n3497 dvss.n527 539.294
R8656 dvss.n3497 dvss.n518 539.294
R8657 dvss.n518 dvss.n510 539.294
R8658 dvss.n3513 dvss.n510 539.294
R8659 dvss.n3563 dvss.n3513 539.294
R8660 dvss.n3518 dvss.n3517 539.294
R8661 dvss.n3568 dvss.n3567 539.294
R8662 dvss.n3568 dvss.n3527 539.294
R8663 dvss.n3528 dvss.n3527 539.294
R8664 dvss.n3575 dvss.n3528 539.294
R8665 dvss.n3576 dvss.n3575 539.294
R8666 dvss.n3576 dvss.n3538 539.294
R8667 dvss.n3539 dvss.n3538 539.294
R8668 dvss.n3545 dvss.n3539 539.294
R8669 dvss.n3545 dvss.n3544 539.294
R8670 dvss.n3544 dvss.n371 539.294
R8671 dvss.n377 dvss.n371 539.294
R8672 dvss.n447 dvss.n377 539.294
R8673 dvss.n449 dvss.n447 539.294
R8674 dvss.n449 dvss.n443 539.294
R8675 dvss.n458 dvss.n443 539.294
R8676 dvss.n458 dvss.n439 539.294
R8677 dvss.n439 dvss.n390 539.294
R8678 dvss.n391 dvss.n390 539.294
R8679 dvss.n430 dvss.n391 539.294
R8680 dvss.n397 dvss.n396 539.294
R8681 dvss.n435 dvss.n434 539.294
R8682 dvss.n435 dvss.n406 539.294
R8683 dvss.n407 dvss.n406 539.294
R8684 dvss.n425 dvss.n407 539.294
R8685 dvss.n426 dvss.n425 539.294
R8686 dvss.n426 dvss.n417 539.294
R8687 dvss.n418 dvss.n417 539.294
R8688 dvss.n3838 dvss.n418 539.294
R8689 dvss.n3840 dvss.n3838 539.294
R8690 dvss.n3840 dvss.n346 539.294
R8691 dvss.n3939 dvss.n346 539.294
R8692 dvss.n3940 dvss.n3939 539.294
R8693 dvss.n3940 dvss.n341 539.294
R8694 dvss.n341 dvss.n330 539.294
R8695 dvss.n3967 dvss.n330 539.294
R8696 dvss.n3968 dvss.n3967 539.294
R8697 dvss.n3968 dvss.n321 539.294
R8698 dvss.n321 dvss.n315 539.294
R8699 dvss.n3982 dvss.n315 539.294
R8700 dvss.n3983 dvss.n3982 539.294
R8701 dvss.n2888 dvss.n2391 539.294
R8702 dvss.n2394 dvss.n2393 539.294
R8703 dvss.n2397 dvss.n2396 539.294
R8704 dvss.n2399 dvss.n2398 539.294
R8705 dvss.n2402 dvss.n2401 539.294
R8706 dvss.n2408 dvss.n2407 539.294
R8707 dvss.n2410 dvss.n2409 539.294
R8708 dvss.n2418 dvss.n2417 539.294
R8709 dvss.n2420 dvss.n2419 539.294
R8710 dvss.n2422 dvss.n2421 539.294
R8711 dvss.n2428 dvss.n2427 539.294
R8712 dvss.n2431 dvss.n2430 539.294
R8713 dvss.n2433 dvss.n2432 539.294
R8714 dvss.n2436 dvss.n2435 539.294
R8715 dvss.n2441 dvss.n2440 539.294
R8716 dvss.n2443 dvss.n2442 539.294
R8717 dvss.n2447 dvss.n2446 539.294
R8718 dvss.n2450 dvss.n2449 539.294
R8719 dvss.n2452 dvss.n2451 539.294
R8720 dvss.n2455 dvss.n2454 539.294
R8721 dvss.n2461 dvss.n2460 539.294
R8722 dvss.n2464 dvss.n2463 539.294
R8723 dvss.n2467 dvss.n2466 539.294
R8724 dvss.n2469 dvss.n2468 539.294
R8725 dvss.n2472 dvss.n2471 539.294
R8726 dvss.n2477 dvss.n2476 539.294
R8727 dvss.n2479 dvss.n2478 539.294
R8728 dvss.n2483 dvss.n2482 539.294
R8729 dvss.n2486 dvss.n2485 539.294
R8730 dvss.n2488 dvss.n2487 539.294
R8731 dvss.n2491 dvss.n2490 539.294
R8732 dvss.n2497 dvss.n2496 539.294
R8733 dvss.n2500 dvss.n2499 539.294
R8734 dvss.n2503 dvss.n2502 539.294
R8735 dvss.n2505 dvss.n2504 539.294
R8736 dvss.n2508 dvss.n2507 539.294
R8737 dvss.n2513 dvss.n2512 539.294
R8738 dvss.n2515 dvss.n2514 539.294
R8739 dvss.n2519 dvss.n2518 539.294
R8740 dvss.n2522 dvss.n2521 539.294
R8741 dvss.n2524 dvss.n2523 539.294
R8742 dvss.n2527 dvss.n2526 539.294
R8743 dvss.n2533 dvss.n2532 539.294
R8744 dvss.n2536 dvss.n2535 539.294
R8745 dvss.n2539 dvss.n2538 539.294
R8746 dvss.n2541 dvss.n2540 539.294
R8747 dvss.n2544 dvss.n2543 539.294
R8748 dvss.n2549 dvss.n2548 539.294
R8749 dvss.n2551 dvss.n2550 539.294
R8750 dvss.n2555 dvss.n2554 539.294
R8751 dvss.n2558 dvss.n2557 539.294
R8752 dvss.n2560 dvss.n2559 539.294
R8753 dvss.n2563 dvss.n2562 539.294
R8754 dvss.n2569 dvss.n2568 539.294
R8755 dvss.n2572 dvss.n2571 539.294
R8756 dvss.n2575 dvss.n2574 539.294
R8757 dvss.n2577 dvss.n2576 539.294
R8758 dvss.n2580 dvss.n2579 539.294
R8759 dvss.n2585 dvss.n2584 539.294
R8760 dvss.n2587 dvss.n2586 539.294
R8761 dvss.n2591 dvss.n2590 539.294
R8762 dvss.n2594 dvss.n2593 539.294
R8763 dvss.n2596 dvss.n2595 539.294
R8764 dvss.n2599 dvss.n2598 539.294
R8765 dvss.n2605 dvss.n2604 539.294
R8766 dvss.n2608 dvss.n2607 539.294
R8767 dvss.n2891 dvss.n2324 539.294
R8768 dvss.n2898 dvss.n2321 539.294
R8769 dvss.n2898 dvss.n2319 539.294
R8770 dvss.n2902 dvss.n2319 539.294
R8771 dvss.n2902 dvss.n2316 539.294
R8772 dvss.n2911 dvss.n2316 539.294
R8773 dvss.n2912 dvss.n2911 539.294
R8774 dvss.n2912 dvss.n2313 539.294
R8775 dvss.n2917 dvss.n2313 539.294
R8776 dvss.n2917 dvss.n2306 539.294
R8777 dvss.n2932 dvss.n2306 539.294
R8778 dvss.n2932 dvss.n2305 539.294
R8779 dvss.n2937 dvss.n2305 539.294
R8780 dvss.n2937 dvss.n2302 539.294
R8781 dvss.n2944 dvss.n2302 539.294
R8782 dvss.n2944 dvss.n2300 539.294
R8783 dvss.n2949 dvss.n2300 539.294
R8784 dvss.n2949 dvss.n2296 539.294
R8785 dvss.n2960 dvss.n2296 539.294
R8786 dvss.n2960 dvss.n2295 539.294
R8787 dvss.n2964 dvss.n2295 539.294
R8788 dvss.n2964 dvss.n2292 539.294
R8789 dvss.n2971 dvss.n2292 539.294
R8790 dvss.n2971 dvss.n2290 539.294
R8791 dvss.n2976 dvss.n2290 539.294
R8792 dvss.n2976 dvss.n2210 539.294
R8793 dvss.n2985 dvss.n2210 539.294
R8794 dvss.n2985 dvss.n2211 539.294
R8795 dvss.n2226 dvss.n2211 539.294
R8796 dvss.n2226 dvss.n2220 539.294
R8797 dvss.n2236 dvss.n2220 539.294
R8798 dvss.n2236 dvss.n2218 539.294
R8799 dvss.n2240 dvss.n2218 539.294
R8800 dvss.n2241 dvss.n2240 539.294
R8801 dvss.n2242 dvss.n2241 539.294
R8802 dvss.n2253 dvss.n2242 539.294
R8803 dvss.n2253 dvss.n2244 539.294
R8804 dvss.n2245 dvss.n2244 539.294
R8805 dvss.n2249 dvss.n2245 539.294
R8806 dvss.n2269 dvss.n2249 539.294
R8807 dvss.n2269 dvss.n2250 539.294
R8808 dvss.n2250 dvss.n260 539.294
R8809 dvss.n261 dvss.n260 539.294
R8810 dvss.n2263 dvss.n261 539.294
R8811 dvss.n2263 dvss.n263 539.294
R8812 dvss.n264 dvss.n263 539.294
R8813 dvss.n2259 dvss.n264 539.294
R8814 dvss.n2259 dvss.n266 539.294
R8815 dvss.n267 dvss.n266 539.294
R8816 dvss.n369 dvss.n267 539.294
R8817 dvss.n369 dvss.n368 539.294
R8818 dvss.n368 dvss.n356 539.294
R8819 dvss.n356 dvss.n350 539.294
R8820 dvss.n3900 dvss.n350 539.294
R8821 dvss.n3901 dvss.n3900 539.294
R8822 dvss.n3901 dvss.n273 539.294
R8823 dvss.n274 dvss.n273 539.294
R8824 dvss.n3905 dvss.n274 539.294
R8825 dvss.n3905 dvss.n276 539.294
R8826 dvss.n277 dvss.n276 539.294
R8827 dvss.n3910 dvss.n277 539.294
R8828 dvss.n3911 dvss.n3910 539.294
R8829 dvss.n3911 dvss.n283 539.294
R8830 dvss.n284 dvss.n283 539.294
R8831 dvss.n3915 dvss.n284 539.294
R8832 dvss.n3915 dvss.n286 539.294
R8833 dvss.n287 dvss.n286 539.294
R8834 dvss.n3919 dvss.n287 539.294
R8835 dvss.n3919 dvss.n289 539.294
R8836 dvss.n290 dvss.n289 539.294
R8837 dvss.n3927 dvss.n290 539.294
R8838 dvss.n3927 dvss.n294 539.294
R8839 dvss.n295 dvss.n294 539.294
R8840 dvss.n3923 dvss.n295 539.294
R8841 dvss.n3923 dvss.n298 539.294
R8842 dvss.n299 dvss.n298 539.294
R8843 dvss.n327 dvss.n299 539.294
R8844 dvss.n327 dvss.n301 539.294
R8845 dvss.n302 dvss.n301 539.294
R8846 dvss.n304 dvss.n302 539.294
R8847 dvss.n4057 dvss.n304 539.294
R8848 dvss.n1197 dvss.n1097 533.678
R8849 dvss.n945 dvss.n940 533.678
R8850 dvss.n1233 dvss.n906 510.284
R8851 dvss.n2255 dvss.n2254 498.113
R8852 dvss.n2256 dvss.n2255 498.113
R8853 dvss.n2268 dvss.n2257 498.113
R8854 dvss.n2267 dvss.n2266 498.113
R8855 dvss.n2266 dvss.n2265 498.113
R8856 dvss.n2265 dvss.n2264 498.113
R8857 dvss.n2264 dvss.n2262 498.113
R8858 dvss.n2945 dvss.n2301 498.113
R8859 dvss.n2946 dvss.n2945 498.113
R8860 dvss.n2948 dvss.n2947 498.113
R8861 dvss.n2962 dvss.n2961 498.113
R8862 dvss.n2963 dvss.n2962 498.113
R8863 dvss.n2963 dvss.n2291 498.113
R8864 dvss.n2972 dvss.n2291 498.113
R8865 dvss.n2973 dvss.n2972 498.113
R8866 dvss.n2262 dvss.n2261 493.485
R8867 dvss.n3981 dvss.n306 491.163
R8868 dvss.t546 dvss 446.038
R8869 dvss.t101 dvss 446.038
R8870 dvss.t554 dvss.n2256 441.038
R8871 dvss.t696 dvss.n2946 441.038
R8872 dvss.n3831 dvss.n424 432.788
R8873 dvss.n3577 dvss.n3574 432.788
R8874 dvss.n3445 dvss.n554 432.788
R8875 dvss.n3327 dvss.n3326 432.788
R8876 dvss.n3214 dvss.n675 432.788
R8877 dvss.n1888 dvss.n1857 432.788
R8878 dvss.n1736 dvss.n784 432.788
R8879 dvss.n1413 dvss.n1382 432.788
R8880 dvss.n1261 dvss.n893 432.788
R8881 dvss.n3823 dvss.t135 410.247
R8882 dvss.n3573 dvss.t469 410.247
R8883 dvss.n3442 dvss.t186 410.247
R8884 dvss.n3323 dvss.t16 410.247
R8885 dvss.n3201 dvss.t636 410.247
R8886 dvss.n1880 dvss.t462 410.247
R8887 dvss.n1723 dvss.t679 410.247
R8888 dvss.n1405 dvss.t511 410.247
R8889 dvss.n1248 dvss.t426 410.247
R8890 dvss.t141 dvss.n3832 401.229
R8891 dvss.t475 dvss.n3580 401.229
R8892 dvss.t192 dvss.n3464 401.229
R8893 dvss.t22 dvss.n3348 401.229
R8894 dvss.n676 dvss.t632 401.229
R8895 dvss.t464 dvss.n1889 401.229
R8896 dvss.n785 dvss.t673 401.229
R8897 dvss.t505 dvss.n1414 401.229
R8898 dvss.n894 dvss.t418 401.229
R8899 dvss.n3821 dvss.n428 396.721
R8900 dvss.n3569 dvss.n3561 396.721
R8901 dvss.n573 dvss.n572 396.721
R8902 dvss.n631 dvss.n630 396.721
R8903 dvss.n3187 dvss.n3186 396.721
R8904 dvss.n1878 dvss.n1861 396.721
R8905 dvss.n1709 dvss.n1708 396.721
R8906 dvss.n1403 dvss.n1386 396.721
R8907 dvss.n1234 dvss.n1233 396.721
R8908 dvss.n2975 dvss.n2973 389.37
R8909 dvss.n2900 dvss.n2899 389.37
R8910 dvss.n943 dvss.n905 380.784
R8911 dvss.n236 dvss.t80 379.31
R8912 dvss.n2254 dvss.n2252 368.271
R8913 dvss.n2936 dvss.n2301 368.271
R8914 dvss.n3981 dvss.n316 358.591
R8915 dvss.n1071 dvss.t233 349.909
R8916 dvss.t246 dvss.n910 349.909
R8917 dvss.n4003 dvss.t693 348.875
R8918 dvss.n2975 dvss.n2974 342.301
R8919 dvss.n2225 dvss.n2224 342.301
R8920 dvss.n2237 dvss.n2219 342.301
R8921 dvss.n2252 dvss.n2251 342.301
R8922 dvss.n2901 dvss.n2900 342.301
R8923 dvss.n2913 dvss.n2314 342.301
R8924 dvss.n2916 dvss.n2914 342.301
R8925 dvss.n2936 dvss.n2935 342.301
R8926 dvss.n3943 dvss.n345 332.075
R8927 dvss.n3971 dvss.n316 332.075
R8928 dvss.n446 dvss.n445 332.075
R8929 dvss.n3812 dvss.n3811 332.075
R8930 dvss.n3492 dvss.n532 332.075
R8931 dvss.n3623 dvss.n511 332.075
R8932 dvss.n3379 dvss.n594 332.075
R8933 dvss.n3405 dvss.n3404 332.075
R8934 dvss.n3260 dvss.n658 332.075
R8935 dvss.n3287 dvss.n3286 332.075
R8936 dvss.n1903 dvss.n1902 332.075
R8937 dvss.n3185 dvss.n689 332.075
R8938 dvss.n1782 dvss.n767 332.075
R8939 dvss.n1965 dvss.n746 332.075
R8940 dvss.n1428 dvss.n1427 332.075
R8941 dvss.n1707 dvss.n798 332.075
R8942 dvss.n1307 dvss.n876 332.075
R8943 dvss.n1490 dvss.n855 332.075
R8944 dvss.t685 dvss.t147 331.955
R8945 dvss.t147 dvss.t481 331.955
R8946 dvss.t235 dvss.t355 327.353
R8947 dvss.t374 dvss.t252 317.724
R8948 dvss.t235 dvss.t98 317.724
R8949 dvss.n2986 dvss.t254 306.646
R8950 dvss.n2315 dvss.t111 306.646
R8951 dvss.n3832 dvss.t139 302.05
R8952 dvss.n3580 dvss.t473 302.05
R8953 dvss.n3464 dvss.t190 302.05
R8954 dvss.n3348 dvss.t20 302.05
R8955 dvss.t634 dvss.n676 302.05
R8956 dvss.n1889 dvss.t458 302.05
R8957 dvss.t675 dvss.n785 302.05
R8958 dvss.n1414 dvss.t509 302.05
R8959 dvss.t424 dvss.n894 302.05
R8960 dvss.n2268 dvss.t556 300.943
R8961 dvss.n2947 dvss.t466 300.943
R8962 dvss.n3932 dvss.t212 297.485
R8963 dvss.n3895 dvss.t123 297.485
R8964 dvss.n2209 dvss.t26 297.485
R8965 dvss.n3365 dvss.t40 297.485
R8966 dvss.n2157 dvss.t299 297.485
R8967 dvss.n1899 dvss.t565 297.485
R8968 dvss.n1608 dvss.t287 297.485
R8969 dvss.n1424 dvss.t590 297.485
R8970 dvss.n1123 dvss.t341 297.485
R8971 dvss.n3823 dvss.t137 293.034
R8972 dvss.t471 dvss.n3573 293.034
R8973 dvss.n3442 dvss.t188 293.034
R8974 dvss.n3323 dvss.t18 293.034
R8975 dvss.n3201 dvss.t638 293.034
R8976 dvss.n1880 dvss.t460 293.034
R8977 dvss.n1723 dvss.t677 293.034
R8978 dvss.n1405 dvss.t507 293.034
R8979 dvss.n1248 dvss.t420 293.034
R8980 dvss.n2238 dvss.t256 292.384
R8981 dvss.t113 dvss.n2915 292.384
R8982 dvss.t688 dvss.t384 284.077
R8983 dvss.n3966 dvss.t214 283.649
R8984 dvss.n457 dvss.t133 283.649
R8985 dvss.n3498 dvss.t28 283.649
R8986 dvss.t42 dvss.n3383 283.649
R8987 dvss.n3267 dvss.t295 283.649
R8988 dvss.n1910 dvss.t569 283.649
R8989 dvss.n1788 dvss.t279 283.649
R8990 dvss.n1435 dvss.t586 283.649
R8991 dvss.n1313 dvss.t337 283.649
R8992 dvss.n4135 dvss.t106 283.474
R8993 dvss.n152 dvss.t167 282.327
R8994 dvss.n255 dvss.t304 282.327
R8995 dvss.n97 dvss.t450 282.327
R8996 dvss.n219 dvss.t553 282.327
R8997 dvss.t602 dvss.t624 281.707
R8998 dvss.t626 dvss.t602 281.707
R8999 dvss.t616 dvss.t626 281.707
R9000 dvss.t628 dvss.t616 281.707
R9001 dvss.t608 dvss.t628 281.707
R9002 dvss.t622 dvss.t608 281.707
R9003 dvss.t612 dvss.t622 281.707
R9004 dvss.t598 dvss.t612 281.707
R9005 dvss.t614 dvss.t598 281.707
R9006 dvss.t600 dvss.t614 281.707
R9007 dvss.t604 dvss.t600 281.707
R9008 dvss.t618 dvss.t604 281.707
R9009 dvss.t620 dvss.t606 281.707
R9010 dvss.t610 dvss.t620 281.707
R9011 dvss.t550 dvss.t546 281.707
R9012 dvss.t548 dvss.t550 281.707
R9013 dvss.t552 dvss.t548 281.707
R9014 dvss.t103 dvss.t101 281.707
R9015 dvss.t107 dvss.t103 281.707
R9016 dvss.t105 dvss.t107 281.707
R9017 dvss.n145 dvss.t163 281.13
R9018 dvss.n248 dvss.t516 281.13
R9019 dvss.n94 dvss.t454 281.13
R9020 dvss.n216 dvss.t547 281.13
R9021 dvss.n4141 dvss.t102 281.13
R9022 dvss.n3812 dvss.n428 276.731
R9023 dvss.n3561 dvss.n511 276.731
R9024 dvss.n3405 dvss.n573 276.731
R9025 dvss.n3287 dvss.n631 276.731
R9026 dvss.n3186 dvss.n3185 276.731
R9027 dvss.n1861 dvss.n746 276.731
R9028 dvss.n1708 dvss.n1707 276.731
R9029 dvss.n1386 dvss.n855 276.731
R9030 dvss.n2261 dvss.n2260 275.899
R9031 dvss.n2260 dvss.n2258 275.899
R9032 dvss.n370 dvss.n353 275.899
R9033 dvss.n3903 dvss.n3902 275.899
R9034 dvss.n3904 dvss.n3903 275.899
R9035 dvss.n3906 dvss.n3904 275.899
R9036 dvss.n3907 dvss.n3906 275.899
R9037 dvss.n3908 dvss.n3907 275.899
R9038 dvss.n3912 dvss.n3909 275.899
R9039 dvss.n3914 dvss.n3913 275.899
R9040 dvss.n3916 dvss.n3914 275.899
R9041 dvss.n3917 dvss.n3916 275.899
R9042 dvss.n3918 dvss.n3917 275.899
R9043 dvss.n3920 dvss.n3918 275.899
R9044 dvss.n3921 dvss.n3920 275.899
R9045 dvss.n3922 dvss.n3921 275.899
R9046 dvss.n3930 dvss.n3929 275.899
R9047 dvss.n328 dvss.n326 275.899
R9048 dvss.n326 dvss.n325 275.899
R9049 dvss.n325 dvss.n305 275.899
R9050 dvss.n4056 dvss.n305 275.899
R9051 dvss.n234 dvss.t618 271.647
R9052 dvss.n58 dvss.n44 270.307
R9053 dvss.n56 dvss.n44 270.307
R9054 dvss.n58 dvss.n57 270.307
R9055 dvss.n57 dvss.n56 270.307
R9056 dvss.t264 dvss.n2238 263.858
R9057 dvss.n2915 dvss.t119 263.858
R9058 dvss dvss.t610 261.586
R9059 dvss.t428 dvss.n3821 261.476
R9060 dvss.t536 dvss.n3569 261.476
R9061 dvss.n572 dvss.t435 261.476
R9062 dvss.n630 dvss.t594 261.476
R9063 dvss.n3187 dvss.t172 261.476
R9064 dvss.t121 dvss.n1878 261.476
R9065 dvss.n1709 dvss.t732 261.476
R9066 dvss.t14 dvss.n1403 261.476
R9067 dvss.n1234 dvss.t12 261.476
R9068 dvss.n2239 dvss.n508 256.726
R9069 dvss.n2934 dvss.n2933 256.726
R9070 dvss.n3966 dvss.t210 255.976
R9071 dvss.n457 dvss.t129 255.976
R9072 dvss.n3498 dvss.t36 255.976
R9073 dvss.n3383 dvss.t48 255.976
R9074 dvss.n3267 dvss.t291 255.976
R9075 dvss.n1910 dvss.t567 255.976
R9076 dvss.n1788 dvss.t281 255.976
R9077 dvss.n1435 dvss.t584 255.976
R9078 dvss.n1313 dvss.t335 255.976
R9079 dvss.n1231 dvss.n1057 255.845
R9080 dvss.n1225 dvss.n1057 255.845
R9081 dvss.n1225 dvss.n1224 255.845
R9082 dvss.n1224 dvss.n1223 255.845
R9083 dvss.n1223 dvss.n1063 255.845
R9084 dvss.n1217 dvss.n1063 255.845
R9085 dvss.n1217 dvss.n1216 255.845
R9086 dvss.n1208 dvss.n1082 255.845
R9087 dvss.n1208 dvss.n1207 255.845
R9088 dvss.n1200 dvss.n1095 255.845
R9089 dvss.n1200 dvss.n1199 255.845
R9090 dvss.n1192 dvss.n1096 255.845
R9091 dvss.n1198 dvss.n1096 253.18
R9092 dvss.n1192 dvss.n1191 252.209
R9093 dvss.t145 dvss.t682 252.159
R9094 dvss.t682 dvss.t656 252.159
R9095 dvss.t656 dvss.t685 252.159
R9096 dvss.n3723 dvss.n3722 251.879
R9097 dvss.n3728 dvss.n3727 251.879
R9098 dvss.n3731 dvss.n3730 251.879
R9099 dvss.n3746 dvss.n3745 251.879
R9100 dvss.n3747 dvss.n3746 251.879
R9101 dvss.n3748 dvss.n3747 251.879
R9102 dvss.n3753 dvss.n3752 251.879
R9103 dvss.n3754 dvss.n3753 251.879
R9104 dvss.n4053 dvss.n308 251.879
R9105 dvss.n3649 dvss.n3648 251.879
R9106 dvss.n3663 dvss.n490 251.879
R9107 dvss.n3666 dvss.n3665 251.879
R9108 dvss.n3679 dvss.n3678 251.879
R9109 dvss.n3681 dvss.n3679 251.879
R9110 dvss.n3681 dvss.n3680 251.879
R9111 dvss.n3695 dvss.n3694 251.879
R9112 dvss.n3695 dvss.n465 251.879
R9113 dvss.n3808 dvss.n466 251.879
R9114 dvss.n2203 dvss.n2202 251.879
R9115 dvss.n2207 dvss.n2206 251.879
R9116 dvss.n2989 dvss.n2988 251.879
R9117 dvss.n2992 dvss.n2991 251.879
R9118 dvss.n2993 dvss.n2992 251.879
R9119 dvss.n2994 dvss.n2993 251.879
R9120 dvss.n2999 dvss.n2998 251.879
R9121 dvss.n2999 dvss.n507 251.879
R9122 dvss.n3627 dvss.n3626 251.879
R9123 dvss.n2178 dvss.n2177 251.879
R9124 dvss.n2182 dvss.n2181 251.879
R9125 dvss.n2185 dvss.n2184 251.879
R9126 dvss.n2188 dvss.n2187 251.879
R9127 dvss.n2189 dvss.n2188 251.879
R9128 dvss.n2190 dvss.n2189 251.879
R9129 dvss.n2195 dvss.n2194 251.879
R9130 dvss.n2197 dvss.n2195 251.879
R9131 dvss.n2200 dvss.n2199 251.879
R9132 dvss.n2150 dvss.n2149 251.879
R9133 dvss.n2155 dvss.n2154 251.879
R9134 dvss.n2160 dvss.n2159 251.879
R9135 dvss.n2163 dvss.n2162 251.879
R9136 dvss.n2164 dvss.n2163 251.879
R9137 dvss.n2165 dvss.n2164 251.879
R9138 dvss.n2170 dvss.n2169 251.879
R9139 dvss.n2172 dvss.n2170 251.879
R9140 dvss.n2175 dvss.n2174 251.879
R9141 dvss.n1991 dvss.n1990 251.879
R9142 dvss.n2005 dvss.n726 251.879
R9143 dvss.n2008 dvss.n2007 251.879
R9144 dvss.n2021 dvss.n2020 251.879
R9145 dvss.n2023 dvss.n2021 251.879
R9146 dvss.n2023 dvss.n2022 251.879
R9147 dvss.n2037 dvss.n2036 251.879
R9148 dvss.n2037 dvss.n701 251.879
R9149 dvss.n3151 dvss.n702 251.879
R9150 dvss.n1601 dvss.n1600 251.879
R9151 dvss.n1606 dvss.n1605 251.879
R9152 dvss.n1611 dvss.n1610 251.879
R9153 dvss.n1614 dvss.n1613 251.879
R9154 dvss.n1615 dvss.n1614 251.879
R9155 dvss.n1616 dvss.n1615 251.879
R9156 dvss.n1621 dvss.n1620 251.879
R9157 dvss.n1621 dvss.n743 251.879
R9158 dvss.n1969 dvss.n1968 251.879
R9159 dvss.n1516 dvss.n1515 251.879
R9160 dvss.n1530 dvss.n835 251.879
R9161 dvss.n1533 dvss.n1532 251.879
R9162 dvss.n1546 dvss.n1545 251.879
R9163 dvss.n1548 dvss.n1546 251.879
R9164 dvss.n1548 dvss.n1547 251.879
R9165 dvss.n1562 dvss.n1561 251.879
R9166 dvss.n1562 dvss.n810 251.879
R9167 dvss.n1673 dvss.n811 251.879
R9168 dvss.n1191 dvss.n1190 251.879
R9169 dvss.n1184 dvss.n1183 251.879
R9170 dvss.n1176 dvss.n1122 251.879
R9171 dvss.n1175 dvss.n1174 251.879
R9172 dvss.n1174 dvss.n1125 251.879
R9173 dvss.n1168 dvss.n1125 251.879
R9174 dvss.n1166 dvss.n1150 251.879
R9175 dvss.n1150 dvss.n852 251.879
R9176 dvss.n1494 dvss.n1493 251.879
R9177 dvss dvss.t552 251.524
R9178 dvss dvss.t105 251.524
R9179 dvss.n3970 dvss.n3969 249.058
R9180 dvss.n3810 dvss.n464 249.058
R9181 dvss.n3624 dvss.n509 249.058
R9182 dvss.n3382 dvss.n576 249.058
R9183 dvss.n3266 dvss.n638 249.058
R9184 dvss.n3154 dvss.n3153 249.058
R9185 dvss.n1966 dvss.n744 249.058
R9186 dvss.n1676 dvss.n1675 249.058
R9187 dvss.n1491 dvss.n853 249.058
R9188 dvss.n1206 dvss.t277 247.851
R9189 dvss.t174 dvss.n355 247.16
R9190 dvss.t665 dvss.n3928 247.16
R9191 dvss.n1023 dvss.t237 245.276
R9192 dvss.n2414 dvss.t249 245.276
R9193 dvss.t227 dvss.n3908 244.286
R9194 dvss.n133 dvss.t729 243.903
R9195 dvss.n174 dvss.t400 240.701
R9196 dvss.n1082 dvss.t268 239.856
R9197 dvss.t231 dvss.n1198 237.19
R9198 dvss.n3998 dvss.t681 236.975
R9199 dvss.n4000 dvss.t684 236.975
R9200 dvss.n48 dvss.t690 236.149
R9201 dvss.n3722 dvss.n3721 230.888
R9202 dvss.n3648 dvss.n498 230.888
R9203 dvss.n2202 dvss.n2201 230.888
R9204 dvss.n2177 dvss.n2176 230.888
R9205 dvss.n2149 dvss.n2148 230.888
R9206 dvss.n1990 dvss.n734 230.888
R9207 dvss.n1600 dvss.n1599 230.888
R9208 dvss.n1515 dvss.n843 230.888
R9209 dvss.n3726 dvss.t10 226.6
R9210 dvss.n3650 dvss.t359 226.6
R9211 dvss.n2205 dvss.t321 226.6
R9212 dvss.n2180 dvss.t52 226.6
R9213 dvss.n2153 dvss.t443 226.6
R9214 dvss.n1992 dvss.t317 226.6
R9215 dvss.n1604 dvss.t648 226.6
R9216 dvss.n1517 dvss.t349 226.6
R9217 dvss.n1115 dvss.t155 226.6
R9218 dvss.n3990 dvss.t687 223.559
R9219 dvss.t6 dvss.n3729 221.619
R9220 dvss.t365 dvss.n3664 221.619
R9221 dvss.t327 dvss.n2208 221.619
R9222 dvss.t58 dvss.n2183 221.619
R9223 dvss.t439 dvss.n2156 221.619
R9224 dvss.t319 dvss.n2006 221.619
R9225 dvss.t642 dvss.n1607 221.619
R9226 dvss.t353 dvss.n1531 221.619
R9227 dvss.n1182 dvss.t157 221.619
R9228 dvss.n3926 dvss.n3925 220.345
R9229 dvss.t383 dvss.t688 218.643
R9230 dvss.n3833 dvss.n422 217.097
R9231 dvss.n3582 dvss.n3581 217.097
R9232 dvss.n3466 dvss.n3465 217.097
R9233 dvss.n3350 dvss.n3349 217.097
R9234 dvss.n3234 dvss.n3233 217.097
R9235 dvss.n1890 dvss.n1855 217.097
R9236 dvss.n1756 dvss.n1755 217.097
R9237 dvss.n1415 dvss.n1380 217.097
R9238 dvss.n1281 dvss.n1280 217.097
R9239 dvss.n1233 dvss.n907 212.969
R9240 dvss.n1233 dvss.n908 212.969
R9241 dvss.n2987 dvss.n2986 210.374
R9242 dvss.n2315 dvss.n600 210.374
R9243 dvss.n4054 dvss.n4053 209.899
R9244 dvss.n3721 dvss.n466 209.899
R9245 dvss.n3626 dvss.n498 209.899
R9246 dvss.n2201 dvss.n2200 209.899
R9247 dvss.n2176 dvss.n2175 209.899
R9248 dvss.n2148 dvss.n702 209.899
R9249 dvss.n1968 dvss.n734 209.899
R9250 dvss.n1599 dvss.n811 209.899
R9251 dvss.n1493 dvss.n843 209.899
R9252 dvss.n4139 dvss.n3 207.213
R9253 dvss.n222 dvss.n218 207.213
R9254 dvss.n150 dvss.n99 207.213
R9255 dvss.n114 dvss.n113 207.213
R9256 dvss.n116 dvss.n115 207.213
R9257 dvss.n122 dvss.n110 207.213
R9258 dvss.n125 dvss.n124 207.213
R9259 dvss.n131 dvss.n107 207.213
R9260 dvss.n105 dvss.n104 207.213
R9261 dvss.n139 dvss.n103 207.213
R9262 dvss.n253 dvss.n7 207.213
R9263 dvss.n22 dvss.n21 207.213
R9264 dvss.n24 dvss.n23 207.213
R9265 dvss.n30 dvss.n18 207.213
R9266 dvss.n33 dvss.n32 207.213
R9267 dvss.n39 dvss.n15 207.213
R9268 dvss.n13 dvss.n12 207.213
R9269 dvss.n242 dvss.n11 207.213
R9270 dvss.n158 dvss.n96 207.213
R9271 dvss.n71 dvss.n70 207.213
R9272 dvss.n75 dvss.n69 207.213
R9273 dvss.n78 dvss.n77 207.213
R9274 dvss.n84 dvss.n66 207.213
R9275 dvss.n87 dvss.n86 207.213
R9276 dvss.n64 dvss.n63 207.213
R9277 dvss.n168 dvss.n92 207.213
R9278 dvss.n191 dvss.n190 207.213
R9279 dvss.n193 dvss.n192 207.213
R9280 dvss.n199 dvss.n187 207.213
R9281 dvss.n202 dvss.n201 207.213
R9282 dvss.n208 dvss.n184 207.213
R9283 dvss.n211 dvss.n210 207.213
R9284 dvss.n232 dvss.n181 207.213
R9285 dvss.n3898 dvss.n3897 204.279
R9286 dvss.n3932 dvss.n3931 204.089
R9287 dvss.n3896 dvss.n3895 204.089
R9288 dvss.n2987 dvss.n2209 204.089
R9289 dvss.n3365 dvss.n600 204.089
R9290 dvss.n2158 dvss.n2157 204.089
R9291 dvss.n1899 dvss.n1898 204.089
R9292 dvss.n1609 dvss.n1608 204.089
R9293 dvss.n1424 dvss.n1423 204.089
R9294 dvss.n1124 dvss.n1123 204.089
R9295 dvss.t486 dvss.t694 202.685
R9296 dvss.t178 dvss.n355 201.177
R9297 dvss.n3928 dvss.t661 201.177
R9298 dvss.n1598 dvss.n1597 200.215
R9299 dvss.n1598 dvss.n1596 200.215
R9300 dvss.n1979 dvss.n1978 200.215
R9301 dvss.n1980 dvss.n1979 200.215
R9302 dvss.n2147 dvss.n2146 200.215
R9303 dvss.n2147 dvss.n2145 200.215
R9304 dvss.n2142 dvss.n2141 200.215
R9305 dvss.n2142 dvss.n2139 200.215
R9306 dvss.n2136 dvss.n2135 200.215
R9307 dvss.n2136 dvss.n2133 200.215
R9308 dvss.n3637 dvss.n3636 200.215
R9309 dvss.n3638 dvss.n3637 200.215
R9310 dvss.n3720 dvss.n3719 200.215
R9311 dvss.n3720 dvss.n3718 200.215
R9312 dvss.n1504 dvss.n1503 200.215
R9313 dvss.n1505 dvss.n1504 200.215
R9314 dvss.n1398 dvss.n1397 200.215
R9315 dvss.n1399 dvss.n1398 200.215
R9316 dvss.n1693 dvss.n797 200.215
R9317 dvss.n1696 dvss.n797 200.215
R9318 dvss.n1873 dvss.n1872 200.215
R9319 dvss.n1874 dvss.n1873 200.215
R9320 dvss.n3171 dvss.n688 200.215
R9321 dvss.n3174 dvss.n688 200.215
R9322 dvss.n3306 dvss.n3305 200.215
R9323 dvss.n3307 dvss.n3306 200.215
R9324 dvss.n3409 dvss.n3408 200.215
R9325 dvss.n3410 dvss.n3409 200.215
R9326 dvss.n3560 dvss.n3559 200.215
R9327 dvss.n3560 dvss.n3555 200.215
R9328 dvss.n3816 dvss.n3815 200.215
R9329 dvss.n3817 dvss.n3816 200.215
R9330 dvss.n1015 dvss.n906 200.215
R9331 dvss.n938 dvss.n906 200.215
R9332 dvss.n944 dvss.n943 200.215
R9333 dvss.n943 dvss.n942 200.215
R9334 dvss.n1390 dvss.n1389 200.215
R9335 dvss.n1391 dvss.n1390 200.215
R9336 dvss.n1689 dvss.n1688 200.215
R9337 dvss.n1688 dvss.n1687 200.215
R9338 dvss.n1865 dvss.n1864 200.215
R9339 dvss.n1866 dvss.n1865 200.215
R9340 dvss.n3167 dvss.n3166 200.215
R9341 dvss.n3166 dvss.n3165 200.215
R9342 dvss.n3294 dvss.n3293 200.215
R9343 dvss.n3295 dvss.n3294 200.215
R9344 dvss.n3419 dvss.n3418 200.215
R9345 dvss.n3420 dvss.n3419 200.215
R9346 dvss.n3565 dvss.n3564 200.215
R9347 dvss.n3566 dvss.n3565 200.215
R9348 dvss.n432 dvss.n431 200.215
R9349 dvss.n433 dvss.n432 200.215
R9350 dvss.n1051 dvss.n908 200.215
R9351 dvss.n1044 dvss.n908 200.215
R9352 dvss.n1042 dvss.n908 200.215
R9353 dvss.n1036 dvss.n908 200.215
R9354 dvss.n1034 dvss.n908 200.215
R9355 dvss.n967 dvss.n907 200.215
R9356 dvss.n977 dvss.n907 200.215
R9357 dvss.n979 dvss.n907 200.215
R9358 dvss.n992 dvss.n907 200.215
R9359 dvss.n994 dvss.n907 200.215
R9360 dvss.n1232 dvss.n1056 200.215
R9361 dvss.n964 dvss.n912 200.215
R9362 dvss.n2889 dvss.n2325 200.215
R9363 dvss.n2889 dvss.n2326 200.215
R9364 dvss.n2889 dvss.n2327 200.215
R9365 dvss.n2889 dvss.n2328 200.215
R9366 dvss.n2889 dvss.n2329 200.215
R9367 dvss.n2889 dvss.n2330 200.215
R9368 dvss.n2889 dvss.n2331 200.215
R9369 dvss.n2889 dvss.n2332 200.215
R9370 dvss.n2889 dvss.n2333 200.215
R9371 dvss.n2889 dvss.n2334 200.215
R9372 dvss.n2889 dvss.n2335 200.215
R9373 dvss.n2889 dvss.n2336 200.215
R9374 dvss.n2889 dvss.n2337 200.215
R9375 dvss.n2889 dvss.n2338 200.215
R9376 dvss.n2889 dvss.n2339 200.215
R9377 dvss.n2889 dvss.n2340 200.215
R9378 dvss.n2889 dvss.n2341 200.215
R9379 dvss.n2889 dvss.n2342 200.215
R9380 dvss.n2889 dvss.n2343 200.215
R9381 dvss.n2889 dvss.n2344 200.215
R9382 dvss.n2889 dvss.n2345 200.215
R9383 dvss.n2889 dvss.n2346 200.215
R9384 dvss.n2889 dvss.n2347 200.215
R9385 dvss.n2889 dvss.n2348 200.215
R9386 dvss.n2889 dvss.n2349 200.215
R9387 dvss.n2889 dvss.n2350 200.215
R9388 dvss.n2889 dvss.n2351 200.215
R9389 dvss.n2889 dvss.n2352 200.215
R9390 dvss.n2889 dvss.n2353 200.215
R9391 dvss.n2889 dvss.n2354 200.215
R9392 dvss.n2889 dvss.n2355 200.215
R9393 dvss.n2889 dvss.n2356 200.215
R9394 dvss.n2889 dvss.n2357 200.215
R9395 dvss.n2889 dvss.n2358 200.215
R9396 dvss.n2889 dvss.n2359 200.215
R9397 dvss.n2889 dvss.n2360 200.215
R9398 dvss.n2889 dvss.n2361 200.215
R9399 dvss.n2889 dvss.n2362 200.215
R9400 dvss.n2889 dvss.n2363 200.215
R9401 dvss.n2889 dvss.n2364 200.215
R9402 dvss.n2889 dvss.n2365 200.215
R9403 dvss.n2889 dvss.n2366 200.215
R9404 dvss.n2889 dvss.n2367 200.215
R9405 dvss.n2889 dvss.n2368 200.215
R9406 dvss.n2889 dvss.n2369 200.215
R9407 dvss.n2889 dvss.n2370 200.215
R9408 dvss.n2889 dvss.n2371 200.215
R9409 dvss.n2889 dvss.n2372 200.215
R9410 dvss.n2889 dvss.n2373 200.215
R9411 dvss.n2889 dvss.n2374 200.215
R9412 dvss.n2889 dvss.n2375 200.215
R9413 dvss.n2889 dvss.n2376 200.215
R9414 dvss.n2889 dvss.n2377 200.215
R9415 dvss.n2889 dvss.n2378 200.215
R9416 dvss.n2889 dvss.n2379 200.215
R9417 dvss.n2889 dvss.n2380 200.215
R9418 dvss.n2889 dvss.n2381 200.215
R9419 dvss.n2889 dvss.n2382 200.215
R9420 dvss.n2889 dvss.n2383 200.215
R9421 dvss.n2889 dvss.n2384 200.215
R9422 dvss.n2889 dvss.n2385 200.215
R9423 dvss.n2889 dvss.n2386 200.215
R9424 dvss.n2889 dvss.n2387 200.215
R9425 dvss.n2889 dvss.n2388 200.215
R9426 dvss.n2889 dvss.n2389 200.215
R9427 dvss.n2889 dvss.n2390 200.215
R9428 dvss.n2890 dvss.n2889 200.215
R9429 dvss.t556 dvss.n2267 197.171
R9430 dvss.n2961 dvss.t466 197.171
R9431 dvss.n4010 dvss.t486 194.704
R9432 dvss.n3754 dvss.n329 188.91
R9433 dvss.n3809 dvss.n465 188.91
R9434 dvss.n3625 dvss.n507 188.91
R9435 dvss.n2198 dvss.n2197 188.91
R9436 dvss.n2173 dvss.n2172 188.91
R9437 dvss.n3152 dvss.n701 188.91
R9438 dvss.n1967 dvss.n743 188.91
R9439 dvss.n1674 dvss.n810 188.91
R9440 dvss.n1492 dvss.n852 188.91
R9441 dvss.t667 dvss.n3924 188.212
R9442 dvss.n3899 dvss.t184 188.212
R9443 dvss.n1022 dvss.n1021 185
R9444 dvss.n2413 dvss.n2412 185
R9445 dvss.n1503 dvss.n1502 184.572
R9446 dvss.n1506 dvss.n1505 184.572
R9447 dvss.n1597 dvss.n1567 184.572
R9448 dvss.n1596 dvss.n1595 184.572
R9449 dvss.n1978 dvss.n1977 184.572
R9450 dvss.n1981 dvss.n1980 184.572
R9451 dvss.n2146 dvss.n2042 184.572
R9452 dvss.n2145 dvss.n2144 184.572
R9453 dvss.n2141 dvss.n2140 184.572
R9454 dvss.n2139 dvss.n2075 184.572
R9455 dvss.n2135 dvss.n2134 184.572
R9456 dvss.n2133 dvss.n2106 184.572
R9457 dvss.n3636 dvss.n3635 184.572
R9458 dvss.n3639 dvss.n3638 184.572
R9459 dvss.n3719 dvss.n3700 184.572
R9460 dvss.n3718 dvss.n3717 184.572
R9461 dvss.n310 dvss.n307 184.572
R9462 dvss.n1597 dvss.n1568 184.572
R9463 dvss.n1596 dvss.n1570 184.572
R9464 dvss.n1978 dvss.n738 184.572
R9465 dvss.n1980 dvss.n735 184.572
R9466 dvss.n2146 dvss.n2043 184.572
R9467 dvss.n2145 dvss.n2045 184.572
R9468 dvss.n2141 dvss.n2074 184.572
R9469 dvss.n2139 dvss.n2138 184.572
R9470 dvss.n2135 dvss.n2105 184.572
R9471 dvss.n2133 dvss.n2132 184.572
R9472 dvss.n3636 dvss.n502 184.572
R9473 dvss.n3638 dvss.n499 184.572
R9474 dvss.n3719 dvss.n3701 184.572
R9475 dvss.n3718 dvss.n3703 184.572
R9476 dvss.n1503 dvss.n847 184.572
R9477 dvss.n1505 dvss.n844 184.572
R9478 dvss.n967 dvss.n966 184.572
R9479 dvss.n977 dvss.n976 184.572
R9480 dvss.n980 dvss.n979 184.572
R9481 dvss.n992 dvss.n991 184.572
R9482 dvss.n995 dvss.n994 184.572
R9483 dvss.n1015 dvss.n1014 184.572
R9484 dvss.n950 dvss.n938 184.572
R9485 dvss.n1397 dvss.n1396 184.572
R9486 dvss.n1400 dvss.n1399 184.572
R9487 dvss.n1693 dvss.n801 184.572
R9488 dvss.n1696 dvss.n1695 184.572
R9489 dvss.n1872 dvss.n1871 184.572
R9490 dvss.n1875 dvss.n1874 184.572
R9491 dvss.n3171 dvss.n692 184.572
R9492 dvss.n3174 dvss.n3173 184.572
R9493 dvss.n3305 dvss.n3304 184.572
R9494 dvss.n3308 dvss.n3307 184.572
R9495 dvss.n3408 dvss.n3407 184.572
R9496 dvss.n3410 dvss.n571 184.572
R9497 dvss.n3559 dvss.n3558 184.572
R9498 dvss.n3555 dvss.n3554 184.572
R9499 dvss.n3815 dvss.n3814 184.572
R9500 dvss.n3818 dvss.n3817 184.572
R9501 dvss.n1397 dvss.n1395 184.572
R9502 dvss.n1399 dvss.n1394 184.572
R9503 dvss.n1694 dvss.n1693 184.572
R9504 dvss.n1697 dvss.n1696 184.572
R9505 dvss.n1872 dvss.n1870 184.572
R9506 dvss.n1874 dvss.n1869 184.572
R9507 dvss.n3172 dvss.n3171 184.572
R9508 dvss.n3175 dvss.n3174 184.572
R9509 dvss.n3305 dvss.n632 184.572
R9510 dvss.n3307 dvss.n629 184.572
R9511 dvss.n3408 dvss.n570 184.572
R9512 dvss.n3411 dvss.n3410 184.572
R9513 dvss.n3559 dvss.n3557 184.572
R9514 dvss.n3556 dvss.n3555 184.572
R9515 dvss.n3815 dvss.n437 184.572
R9516 dvss.n3817 dvss.n436 184.572
R9517 dvss.n1016 dvss.n1015 184.572
R9518 dvss.n938 dvss.n937 184.572
R9519 dvss.n1052 dvss.n1051 184.572
R9520 dvss.n1044 dvss.n918 184.572
R9521 dvss.n1043 dvss.n1042 184.572
R9522 dvss.n1036 dvss.n923 184.572
R9523 dvss.n1035 dvss.n1034 184.572
R9524 dvss.n944 dvss.n941 184.572
R9525 dvss.n942 dvss.n940 184.572
R9526 dvss.n1389 dvss.n1388 184.572
R9527 dvss.n1392 dvss.n1391 184.572
R9528 dvss.n1689 dvss.n1685 184.572
R9529 dvss.n1687 dvss.n795 184.572
R9530 dvss.n1864 dvss.n1863 184.572
R9531 dvss.n1867 dvss.n1866 184.572
R9532 dvss.n3167 dvss.n3163 184.572
R9533 dvss.n3165 dvss.n686 184.572
R9534 dvss.n3293 dvss.n3289 184.572
R9535 dvss.n3295 dvss.n3291 184.572
R9536 dvss.n3418 dvss.n3417 184.572
R9537 dvss.n3421 dvss.n3420 184.572
R9538 dvss.n3564 dvss.n3563 184.572
R9539 dvss.n3567 dvss.n3566 184.572
R9540 dvss.n431 dvss.n430 184.572
R9541 dvss.n434 dvss.n433 184.572
R9542 dvss.n945 dvss.n944 184.572
R9543 dvss.n942 dvss.n904 184.572
R9544 dvss.n1389 dvss.n1332 184.572
R9545 dvss.n1391 dvss.n1333 184.572
R9546 dvss.n1690 dvss.n1689 184.572
R9547 dvss.n1687 dvss.n1686 184.572
R9548 dvss.n1864 dvss.n1807 184.572
R9549 dvss.n1866 dvss.n1808 184.572
R9550 dvss.n3168 dvss.n3167 184.572
R9551 dvss.n3165 dvss.n3164 184.572
R9552 dvss.n3293 dvss.n3290 184.572
R9553 dvss.n3296 dvss.n3295 184.572
R9554 dvss.n3418 dvss.n564 184.572
R9555 dvss.n3420 dvss.n562 184.572
R9556 dvss.n3564 dvss.n3517 184.572
R9557 dvss.n3566 dvss.n3518 184.572
R9558 dvss.n431 dvss.n396 184.572
R9559 dvss.n433 dvss.n397 184.572
R9560 dvss.n1051 dvss.n1050 184.572
R9561 dvss.n1045 dvss.n1044 184.572
R9562 dvss.n1042 dvss.n1041 184.572
R9563 dvss.n1037 dvss.n1036 184.572
R9564 dvss.n1034 dvss.n1033 184.572
R9565 dvss.n968 dvss.n967 184.572
R9566 dvss.n978 dvss.n977 184.572
R9567 dvss.n979 dvss.n955 184.572
R9568 dvss.n993 dvss.n992 184.572
R9569 dvss.n994 dvss.n952 184.572
R9570 dvss.n1056 dvss.n913 184.572
R9571 dvss.n965 dvss.n964 184.572
R9572 dvss.n2391 dvss.n2325 184.572
R9573 dvss.n2394 dvss.n2326 184.572
R9574 dvss.n2397 dvss.n2327 184.572
R9575 dvss.n2399 dvss.n2328 184.572
R9576 dvss.n2402 dvss.n2329 184.572
R9577 dvss.n2408 dvss.n2330 184.572
R9578 dvss.n2410 dvss.n2331 184.572
R9579 dvss.n2418 dvss.n2332 184.572
R9580 dvss.n2420 dvss.n2333 184.572
R9581 dvss.n2422 dvss.n2334 184.572
R9582 dvss.n2428 dvss.n2335 184.572
R9583 dvss.n2431 dvss.n2336 184.572
R9584 dvss.n2433 dvss.n2337 184.572
R9585 dvss.n2436 dvss.n2338 184.572
R9586 dvss.n2441 dvss.n2339 184.572
R9587 dvss.n2443 dvss.n2340 184.572
R9588 dvss.n2447 dvss.n2341 184.572
R9589 dvss.n2450 dvss.n2342 184.572
R9590 dvss.n2452 dvss.n2343 184.572
R9591 dvss.n2455 dvss.n2344 184.572
R9592 dvss.n2461 dvss.n2345 184.572
R9593 dvss.n2464 dvss.n2346 184.572
R9594 dvss.n2467 dvss.n2347 184.572
R9595 dvss.n2469 dvss.n2348 184.572
R9596 dvss.n2472 dvss.n2349 184.572
R9597 dvss.n2477 dvss.n2350 184.572
R9598 dvss.n2479 dvss.n2351 184.572
R9599 dvss.n2483 dvss.n2352 184.572
R9600 dvss.n2486 dvss.n2353 184.572
R9601 dvss.n2488 dvss.n2354 184.572
R9602 dvss.n2491 dvss.n2355 184.572
R9603 dvss.n2497 dvss.n2356 184.572
R9604 dvss.n2500 dvss.n2357 184.572
R9605 dvss.n2503 dvss.n2358 184.572
R9606 dvss.n2505 dvss.n2359 184.572
R9607 dvss.n2508 dvss.n2360 184.572
R9608 dvss.n2513 dvss.n2361 184.572
R9609 dvss.n2515 dvss.n2362 184.572
R9610 dvss.n2519 dvss.n2363 184.572
R9611 dvss.n2522 dvss.n2364 184.572
R9612 dvss.n2524 dvss.n2365 184.572
R9613 dvss.n2527 dvss.n2366 184.572
R9614 dvss.n2533 dvss.n2367 184.572
R9615 dvss.n2536 dvss.n2368 184.572
R9616 dvss.n2539 dvss.n2369 184.572
R9617 dvss.n2541 dvss.n2370 184.572
R9618 dvss.n2544 dvss.n2371 184.572
R9619 dvss.n2549 dvss.n2372 184.572
R9620 dvss.n2551 dvss.n2373 184.572
R9621 dvss.n2555 dvss.n2374 184.572
R9622 dvss.n2558 dvss.n2375 184.572
R9623 dvss.n2560 dvss.n2376 184.572
R9624 dvss.n2563 dvss.n2377 184.572
R9625 dvss.n2569 dvss.n2378 184.572
R9626 dvss.n2572 dvss.n2379 184.572
R9627 dvss.n2575 dvss.n2380 184.572
R9628 dvss.n2577 dvss.n2381 184.572
R9629 dvss.n2580 dvss.n2382 184.572
R9630 dvss.n2585 dvss.n2383 184.572
R9631 dvss.n2587 dvss.n2384 184.572
R9632 dvss.n2591 dvss.n2385 184.572
R9633 dvss.n2594 dvss.n2386 184.572
R9634 dvss.n2596 dvss.n2387 184.572
R9635 dvss.n2599 dvss.n2388 184.572
R9636 dvss.n2605 dvss.n2389 184.572
R9637 dvss.n2608 dvss.n2390 184.572
R9638 dvss.n2891 dvss.n2890 184.572
R9639 dvss.n2393 dvss.n2325 184.572
R9640 dvss.n2396 dvss.n2326 184.572
R9641 dvss.n2398 dvss.n2327 184.572
R9642 dvss.n2401 dvss.n2328 184.572
R9643 dvss.n2407 dvss.n2329 184.572
R9644 dvss.n2409 dvss.n2330 184.572
R9645 dvss.n2417 dvss.n2331 184.572
R9646 dvss.n2419 dvss.n2332 184.572
R9647 dvss.n2421 dvss.n2333 184.572
R9648 dvss.n2427 dvss.n2334 184.572
R9649 dvss.n2430 dvss.n2335 184.572
R9650 dvss.n2432 dvss.n2336 184.572
R9651 dvss.n2435 dvss.n2337 184.572
R9652 dvss.n2440 dvss.n2338 184.572
R9653 dvss.n2442 dvss.n2339 184.572
R9654 dvss.n2446 dvss.n2340 184.572
R9655 dvss.n2449 dvss.n2341 184.572
R9656 dvss.n2451 dvss.n2342 184.572
R9657 dvss.n2454 dvss.n2343 184.572
R9658 dvss.n2460 dvss.n2344 184.572
R9659 dvss.n2463 dvss.n2345 184.572
R9660 dvss.n2466 dvss.n2346 184.572
R9661 dvss.n2468 dvss.n2347 184.572
R9662 dvss.n2471 dvss.n2348 184.572
R9663 dvss.n2476 dvss.n2349 184.572
R9664 dvss.n2478 dvss.n2350 184.572
R9665 dvss.n2482 dvss.n2351 184.572
R9666 dvss.n2485 dvss.n2352 184.572
R9667 dvss.n2487 dvss.n2353 184.572
R9668 dvss.n2490 dvss.n2354 184.572
R9669 dvss.n2496 dvss.n2355 184.572
R9670 dvss.n2499 dvss.n2356 184.572
R9671 dvss.n2502 dvss.n2357 184.572
R9672 dvss.n2504 dvss.n2358 184.572
R9673 dvss.n2507 dvss.n2359 184.572
R9674 dvss.n2512 dvss.n2360 184.572
R9675 dvss.n2514 dvss.n2361 184.572
R9676 dvss.n2518 dvss.n2362 184.572
R9677 dvss.n2521 dvss.n2363 184.572
R9678 dvss.n2523 dvss.n2364 184.572
R9679 dvss.n2526 dvss.n2365 184.572
R9680 dvss.n2532 dvss.n2366 184.572
R9681 dvss.n2535 dvss.n2367 184.572
R9682 dvss.n2538 dvss.n2368 184.572
R9683 dvss.n2540 dvss.n2369 184.572
R9684 dvss.n2543 dvss.n2370 184.572
R9685 dvss.n2548 dvss.n2371 184.572
R9686 dvss.n2550 dvss.n2372 184.572
R9687 dvss.n2554 dvss.n2373 184.572
R9688 dvss.n2557 dvss.n2374 184.572
R9689 dvss.n2559 dvss.n2375 184.572
R9690 dvss.n2562 dvss.n2376 184.572
R9691 dvss.n2568 dvss.n2377 184.572
R9692 dvss.n2571 dvss.n2378 184.572
R9693 dvss.n2574 dvss.n2379 184.572
R9694 dvss.n2576 dvss.n2380 184.572
R9695 dvss.n2579 dvss.n2381 184.572
R9696 dvss.n2584 dvss.n2382 184.572
R9697 dvss.n2586 dvss.n2383 184.572
R9698 dvss.n2590 dvss.n2384 184.572
R9699 dvss.n2593 dvss.n2385 184.572
R9700 dvss.n2595 dvss.n2386 184.572
R9701 dvss.n2598 dvss.n2387 184.572
R9702 dvss.n2604 dvss.n2388 184.572
R9703 dvss.n2607 dvss.n2389 184.572
R9704 dvss.n2390 dvss.n2324 184.572
R9705 dvss.n2890 dvss.n2321 184.572
R9706 dvss.n2225 dvss.t262 178.282
R9707 dvss.t117 dvss.n2913 178.282
R9708 dvss.n3943 dvss.t206 172.957
R9709 dvss.n446 dvss.t131 172.957
R9710 dvss.n3492 dvss.t34 172.957
R9711 dvss.t46 dvss.n3379 172.957
R9712 dvss.n3260 dvss.t297 172.957
R9713 dvss.n1903 dvss.t571 172.957
R9714 dvss.n1782 dvss.t285 172.957
R9715 dvss.n1428 dvss.t588 172.957
R9716 dvss.n1307 dvss.t339 172.957
R9717 dvss.n3822 dvss.t428 171.311
R9718 dvss.n3570 dvss.t536 171.311
R9719 dvss.n3441 dvss.t435 171.311
R9720 dvss.n3322 dvss.t594 171.311
R9721 dvss.n3200 dvss.t172 171.311
R9722 dvss.n1879 dvss.t121 171.311
R9723 dvss.n1722 dvss.t732 171.311
R9724 dvss.n1404 dvss.t14 171.311
R9725 dvss.n1247 dvss.t12 171.311
R9726 dvss.n3924 dvss.t663 169.85
R9727 dvss.n3899 dvss.t180 169.85
R9728 dvss.n3942 dvss.t499 169.498
R9729 dvss.n450 dvss.t495 169.498
R9730 dvss.t519 dvss.n3495 169.498
R9731 dvss.t370 dvss.n3380 169.498
R9732 dvss.t96 dvss.n3263 169.498
R9733 dvss.n1906 dvss.t640 169.498
R9734 dvss.t513 dvss.n1785 169.498
R9735 dvss.n1431 dvss.t432 169.498
R9736 dvss.t490 dvss.n1310 169.498
R9737 dvss.t271 dvss.n1206 167.899
R9738 dvss.n3729 dvss.t4 166.838
R9739 dvss.n3664 dvss.t363 166.838
R9740 dvss.n2208 dvss.t325 166.838
R9741 dvss.n2183 dvss.t56 166.838
R9742 dvss.n2156 dvss.t441 166.838
R9743 dvss.n2006 dvss.t313 166.838
R9744 dvss.n1607 dvss.t644 166.838
R9745 dvss.n1531 dvss.t347 166.838
R9746 dvss.t153 dvss.n1182 166.838
R9747 dvss.t229 dvss.n3912 166.689
R9748 dvss.t262 dvss.n2219 164.019
R9749 dvss.n2914 dvss.t117 164.019
R9750 dvss.t499 dvss.n3941 162.579
R9751 dvss.n456 dvss.t495 162.579
R9752 dvss.n3496 dvss.t519 162.579
R9753 dvss.n3384 dvss.t370 162.579
R9754 dvss.n3264 dvss.t96 162.579
R9755 dvss.n1909 dvss.t640 162.579
R9756 dvss.n1786 dvss.t513 162.579
R9757 dvss.n1434 dvss.t432 162.579
R9758 dvss.n1311 dvss.t490 162.579
R9759 dvss.n3712 dvss 161.882
R9760 dvss.n3657 dvss 161.882
R9761 dvss.n2116 dvss 161.882
R9762 dvss.n2085 dvss 161.882
R9763 dvss.n2054 dvss 161.882
R9764 dvss.n1999 dvss 161.882
R9765 dvss.n1579 dvss 161.882
R9766 dvss.n1524 dvss 161.882
R9767 dvss.n1132 dvss 161.882
R9768 dvss.n3857 dvss 161.882
R9769 dvss.n3601 dvss 161.882
R9770 dvss.n549 dvss 161.882
R9771 dvss.n3333 dvss 161.882
R9772 dvss.n672 dvss 161.882
R9773 dvss.n1943 dvss 161.882
R9774 dvss.n781 dvss 161.882
R9775 dvss.n1468 dvss 161.882
R9776 dvss.n890 dvss 161.882
R9777 dvss.t2 dvss.n3726 161.857
R9778 dvss.n3650 dvss.t361 161.857
R9779 dvss.t323 dvss.n2205 161.857
R9780 dvss.t54 dvss.n2180 161.857
R9781 dvss.t445 dvss.n2153 161.857
R9782 dvss.n1992 dvss.t315 161.857
R9783 dvss.t646 dvss.n1604 161.857
R9784 dvss.n1517 dvss.t345 161.857
R9785 dvss.t149 dvss.n1115 161.857
R9786 dvss.n112 dvss.t708 161.522
R9787 dvss.n72 dvss.t411 161.522
R9788 dvss.n20 dvss.t91 161.47
R9789 dvss.n189 dvss.t625 161.143
R9790 dvss.n1084 dvss.t276 160.064
R9791 dvss.n998 dvss.t380 160.064
R9792 dvss.n1216 dvss.n1215 157.238
R9793 dvss.n3748 dvss.t216 154.8
R9794 dvss.n3680 dvss.t125 154.8
R9795 dvss.n2994 dvss.t30 154.8
R9796 dvss.n2190 dvss.t44 154.8
R9797 dvss.n2165 dvss.t293 154.8
R9798 dvss.n2022 dvss.t563 154.8
R9799 dvss.n1616 dvss.t283 154.8
R9800 dvss.n1547 dvss.t582 154.8
R9801 dvss.n1168 dvss.t333 154.8
R9802 dvss.n1075 dvss.t269 154.305
R9803 dvss.n985 dvss.t502 154.305
R9804 dvss.t694 dvss.t383 153.21
R9805 dvss.n101 dvss.t718 152.838
R9806 dvss.n9 dvss.t69 152.838
R9807 dvss.n93 dvss.t389 152.838
R9808 dvss.n215 dvss.t611 152.838
R9809 dvss.n3839 dvss.t143 148.743
R9810 dvss.n3543 dvss.t477 148.743
R9811 dvss.n3470 dvss.t194 148.743
R9812 dvss.t24 dvss.n608 148.743
R9813 dvss.n3238 dvss.t630 148.743
R9814 dvss.n1897 dvss.t456 148.743
R9815 dvss.n1760 dvss.t671 148.743
R9816 dvss.n1422 dvss.t503 148.743
R9817 dvss.n1285 dvss.t422 148.743
R9818 dvss.n56 dvss.n55 146.25
R9819 dvss.n55 dvss.n54 146.25
R9820 dvss.n59 dvss.n58 146.25
R9821 dvss.n60 dvss.n59 146.25
R9822 dvss.t182 dvss.n353 143.697
R9823 dvss.n3929 dvss.t659 143.697
R9824 dvss.t137 dvss.n424 139.755
R9825 dvss.n3574 dvss.t471 139.755
R9826 dvss.n3445 dvss.t188 139.755
R9827 dvss.n3327 dvss.t18 139.755
R9828 dvss.t638 dvss.n675 139.755
R9829 dvss.t460 dvss.n1857 139.755
R9830 dvss.t677 dvss.n784 139.755
R9831 dvss.t507 dvss.n1382 139.755
R9832 dvss.t420 dvss.n893 139.755
R9833 dvss.n1003 dvss.t234 139.52
R9834 dvss.n2404 dvss.t247 139.52
R9835 dvss.n3731 dvss.t8 139.059
R9836 dvss.n3665 dvss.t367 139.059
R9837 dvss.t329 dvss.n2989 139.059
R9838 dvss.t60 dvss.n2185 139.059
R9839 dvss.t437 dvss.n2160 139.059
R9840 dvss.n2007 dvss.t311 139.059
R9841 dvss.t650 dvss.n1611 139.059
R9842 dvss.n1532 dvss.t351 139.059
R9843 dvss.n1176 dvss.t151 139.059
R9844 dvss.n1084 dvss.t274 137.442
R9845 dvss.n1085 dvss.t272 137.442
R9846 dvss.n998 dvss.t378 137.442
R9847 dvss.n999 dvss.t376 137.442
R9848 dvss.n422 dvss.t143 134.488
R9849 dvss.n3582 dvss.t477 134.488
R9850 dvss.n3466 dvss.t194 134.488
R9851 dvss.n3350 dvss.t24 134.488
R9852 dvss.n3234 dvss.t630 134.488
R9853 dvss.n1855 dvss.t456 134.488
R9854 dvss.n1756 dvss.t671 134.488
R9855 dvss.n1380 dvss.t503 134.488
R9856 dvss.n1281 dvss.t422 134.488
R9857 dvss.t182 dvss.n354 132.202
R9858 dvss.t139 dvss.n3831 130.738
R9859 dvss.n3577 dvss.t473 130.738
R9860 dvss.n554 dvss.t190 130.738
R9861 dvss.n3326 dvss.t20 130.738
R9862 dvss.n3214 dvss.t634 130.738
R9863 dvss.t458 dvss.n1888 130.738
R9864 dvss.n1736 dvss.t675 130.738
R9865 dvss.t509 dvss.n1413 130.738
R9866 dvss.n1261 dvss.t424 130.738
R9867 dvss.t50 dvss.n3751 128.564
R9868 dvss.t497 dvss.n3693 128.564
R9869 dvss.t225 dvss.n2997 128.564
R9870 dvss.t309 dvss.n2193 128.564
R9871 dvss.t524 dvss.n2168 128.564
R9872 dvss.t492 dvss.n2035 128.564
R9873 dvss.t430 dvss.n1619 128.564
R9874 dvss.t521 dvss.n1560 128.564
R9875 dvss.n1167 dvss.t372 128.564
R9876 dvss.t669 dvss.n3942 127.987
R9877 dvss.n450 dvss.t176 127.987
R9878 dvss.n3495 dvss.t258 127.987
R9879 dvss.n3380 dvss.t115 127.987
R9880 dvss.n3263 dvss.t539 127.987
R9881 dvss.n1906 dvss.t575 127.987
R9882 dvss.n1785 dvss.t529 127.987
R9883 dvss.n1431 dvss.t198 127.987
R9884 dvss.n1310 dvss.t239 127.987
R9885 dvss.n3931 dvss.t661 125.389
R9886 dvss.n3896 dvss.t178 125.389
R9887 dvss.n3752 dvss.t50 123.316
R9888 dvss.n3694 dvss.t497 123.316
R9889 dvss.n2998 dvss.t225 123.316
R9890 dvss.n2194 dvss.t309 123.316
R9891 dvss.n2169 dvss.t524 123.316
R9892 dvss.n2036 dvss.t492 123.316
R9893 dvss.n1620 dvss.t430 123.316
R9894 dvss.n1561 dvss.t521 123.316
R9895 dvss.t372 dvss.n1166 123.316
R9896 dvss.n3960 dvss.t211 116.939
R9897 dvss.n3878 dvss.t130 116.939
R9898 dvss.n3509 dvss.t37 116.939
R9899 dvss.n3395 dvss.t49 116.939
R9900 dvss.n3278 dvss.t292 116.939
R9901 dvss.n3159 dvss.t568 116.939
R9902 dvss.n1799 dvss.t282 116.939
R9903 dvss.n1681 dvss.t585 116.939
R9904 dvss.n1324 dvss.t336 116.939
R9905 dvss.n4066 dvss.t664 116.939
R9906 dvss.n4113 dvss.t181 116.939
R9907 dvss.n2286 dvss.t265 116.939
R9908 dvss.n2928 dvss.t120 116.939
R9909 dvss.n2628 dvss.t538 116.939
R9910 dvss.n2675 dvss.t578 116.939
R9911 dvss.n2722 dvss.t528 116.939
R9912 dvss.n2769 dvss.t201 116.939
R9913 dvss.n2816 dvss.t241 116.939
R9914 dvss.n3775 dvss.t9 116.938
R9915 dvss.n3673 dvss.t368 116.938
R9916 dvss.n3018 dvss.t330 116.938
R9917 dvss.n3068 dvss.t61 116.938
R9918 dvss.n3118 dvss.t438 116.938
R9919 dvss.n2015 dvss.t312 116.938
R9920 dvss.n1640 dvss.t651 116.938
R9921 dvss.n1540 dvss.t352 116.938
R9922 dvss.n1143 dvss.t152 116.938
R9923 dvss.n3848 dvss.t144 116.938
R9924 dvss.n3592 dvss.t478 116.938
R9925 dvss.n3475 dvss.t195 116.938
R9926 dvss.n3359 dvss.t25 116.938
R9927 dvss.n3243 dvss.t631 116.938
R9928 dvss.n1934 dvss.t457 116.938
R9929 dvss.n1765 dvss.t672 116.938
R9930 dvss.n1459 dvss.t504 116.938
R9931 dvss.n1290 dvss.t423 116.938
R9932 dvss.n1124 dvss.t200 116.547
R9933 dvss.n1609 dvss.t200 116.547
R9934 dvss.n2158 dvss.t200 116.547
R9935 dvss.n1898 dvss.t200 116.547
R9936 dvss.n1423 dvss.t200 116.547
R9937 dvss dvss.n3739 113.316
R9938 dvss dvss.n475 113.316
R9939 dvss dvss.n2127 113.316
R9940 dvss dvss.n2096 113.316
R9941 dvss dvss.n2065 113.316
R9942 dvss dvss.n711 113.316
R9943 dvss dvss.n1590 113.316
R9944 dvss dvss.n820 113.316
R9945 dvss dvss.n1153 113.316
R9946 dvss dvss.n3948 113.316
R9947 dvss dvss.n381 113.316
R9948 dvss dvss.n3483 113.316
R9949 dvss dvss.n3372 113.316
R9950 dvss dvss.n3251 113.316
R9951 dvss dvss.n1846 113.316
R9952 dvss dvss.n1773 113.316
R9953 dvss dvss.n1371 113.316
R9954 dvss dvss.n1298 113.316
R9955 dvss.n3745 dvss.t8 112.822
R9956 dvss.n3678 dvss.t367 112.822
R9957 dvss.n2991 dvss.t329 112.822
R9958 dvss.n2187 dvss.t60 112.822
R9959 dvss.n2162 dvss.t437 112.822
R9960 dvss.n2020 dvss.t311 112.822
R9961 dvss.n1613 dvss.t650 112.822
R9962 dvss.n1545 dvss.t351 112.822
R9963 dvss.t151 dvss.n1175 112.822
R9964 dvss.n3913 dvss.t229 109.21
R9965 dvss.n2899 dvss.n2320 108.963
R9966 dvss.n1100 dvss.n1098 105.862
R9967 dvss.n1027 dvss.n1020 105.862
R9968 dvss.t659 dvss.n3926 105.582
R9969 dvss.n1215 dvss.n1214 98.6074
R9970 dvss.n3751 dvss.t216 97.0786
R9971 dvss.n3693 dvss.t125 97.0786
R9972 dvss.n2997 dvss.t30 97.0786
R9973 dvss.n2193 dvss.t44 97.0786
R9974 dvss.n2168 dvss.t293 97.0786
R9975 dvss.n2035 dvss.t563 97.0786
R9976 dvss.n1619 dvss.t283 97.0786
R9977 dvss.n1560 dvss.t582 97.0786
R9978 dvss.t333 dvss.n1167 97.0786
R9979 dvss.n2974 dvss.t260 92.7071
R9980 dvss.n2901 dvss.t109 92.7071
R9981 dvss.n402 dvss.n401 90.0716
R9982 dvss.n3523 dvss.n3522 90.0716
R9983 dvss.n3426 dvss.n3425 90.0716
R9984 dvss.n3313 dvss.n3312 90.0716
R9985 dvss.n3194 dvss.n3193 90.0716
R9986 dvss.n1813 dvss.n1812 90.0716
R9987 dvss.n1716 dvss.n1715 90.0716
R9988 dvss.n1338 dvss.n1337 90.0716
R9989 dvss.n1241 dvss.n1240 90.0716
R9990 dvss.n1005 dvss.n1004 90.0716
R9991 dvss.n280 dvss.n279 90.0716
R9992 dvss.n2248 dvss.n2247 90.0716
R9993 dvss.n2954 dvss.n2953 90.0716
R9994 dvss.n2602 dvss.n2601 90.0716
R9995 dvss.n2566 dvss.n2565 90.0716
R9996 dvss.n2530 dvss.n2529 90.0716
R9997 dvss.n2494 dvss.n2493 90.0716
R9998 dvss.n2458 dvss.n2457 90.0716
R9999 dvss.n2425 dvss.n2424 90.0716
R10000 dvss.n2406 dvss.n2405 90.0716
R10001 dvss.n3839 dvss.t208 89.9376
R10002 dvss.n3543 dvss.t127 89.9376
R10003 dvss.n3470 dvss.t32 89.9376
R10004 dvss.n608 dvss.t38 89.9376
R10005 dvss.n3238 dvss.t301 89.9376
R10006 dvss.t573 dvss.n1897 89.9376
R10007 dvss.n1760 dvss.t289 89.9376
R10008 dvss.t592 dvss.n1422 89.9376
R10009 dvss.n1285 dvss.t343 89.9376
R10010 dvss.n1207 dvss.t271 87.9472
R10011 dvss.n2251 dvss.n508 85.5759
R10012 dvss.n2935 dvss.n2934 85.5759
R10013 dvss.n51 dvss.t219 84.171
R10014 dvss.n3971 dvss.n3970 83.0194
R10015 dvss.n3811 dvss.n3810 83.0194
R10016 dvss.n3624 dvss.n3623 83.0194
R10017 dvss.n3404 dvss.n576 83.0194
R10018 dvss.n3286 dvss.n638 83.0194
R10019 dvss.n3153 dvss.n689 83.0194
R10020 dvss.n1966 dvss.n1965 83.0194
R10021 dvss.n1675 dvss.n798 83.0194
R10022 dvss.n1491 dvss.n1490 83.0194
R10023 dvss.n3727 dvss.t2 81.3362
R10024 dvss.n490 dvss.t361 81.3362
R10025 dvss.n2206 dvss.t323 81.3362
R10026 dvss.n2181 dvss.t54 81.3362
R10027 dvss.n2154 dvss.t445 81.3362
R10028 dvss.n726 dvss.t315 81.3362
R10029 dvss.n1605 dvss.t646 81.3362
R10030 dvss.n835 dvss.t345 81.3362
R10031 dvss.n1184 dvss.t149 81.3362
R10032 dvss.n4013 dvss.n4012 79.7974
R10033 dvss.n2239 dvss.t264 78.4446
R10034 dvss.n2933 dvss.t119 78.4446
R10035 dvss.n3959 dvss.n335 76.7239
R10036 dvss.n3960 dvss.n3959 76.7239
R10037 dvss.n3879 dvss.n386 76.7239
R10038 dvss.n3879 dvss.n3878 76.7239
R10039 dvss.n3508 dvss.n520 76.7239
R10040 dvss.n3509 dvss.n3508 76.7239
R10041 dvss.n3394 dvss.n583 76.7239
R10042 dvss.n3395 dvss.n3394 76.7239
R10043 dvss.n3277 dvss.n646 76.7239
R10044 dvss.n3278 dvss.n3277 76.7239
R10045 dvss.n1841 dvss.n697 76.7239
R10046 dvss.n3159 dvss.n697 76.7239
R10047 dvss.n1798 dvss.n755 76.7239
R10048 dvss.n1799 dvss.n1798 76.7239
R10049 dvss.n1366 dvss.n806 76.7239
R10050 dvss.n1681 dvss.n806 76.7239
R10051 dvss.n1323 dvss.n864 76.7239
R10052 dvss.n1324 dvss.n1323 76.7239
R10053 dvss.n4083 dvss.n292 76.7239
R10054 dvss.n4066 dvss.n292 76.7239
R10055 dvss.n4117 dvss.n4114 76.7239
R10056 dvss.n4114 dvss.n4113 76.7239
R10057 dvss.n2981 dvss.n2287 76.7239
R10058 dvss.n2287 dvss.n2286 76.7239
R10059 dvss.n2925 dvss.n2309 76.7239
R10060 dvss.n2928 dvss.n2925 76.7239
R10061 dvss.n2645 dvss.n2582 76.7239
R10062 dvss.n2628 dvss.n2582 76.7239
R10063 dvss.n2692 dvss.n2546 76.7239
R10064 dvss.n2675 dvss.n2546 76.7239
R10065 dvss.n2739 dvss.n2510 76.7239
R10066 dvss.n2722 dvss.n2510 76.7239
R10067 dvss.n2786 dvss.n2474 76.7239
R10068 dvss.n2769 dvss.n2474 76.7239
R10069 dvss.n2833 dvss.n2438 76.7239
R10070 dvss.n2816 dvss.n2438 76.7239
R10071 dvss.n3969 dvss.t210 76.1011
R10072 dvss.n464 dvss.t129 76.1011
R10073 dvss.t36 dvss.n509 76.1011
R10074 dvss.t48 dvss.n3382 76.1011
R10075 dvss.t291 dvss.n3266 76.1011
R10076 dvss.n3154 dvss.t567 76.1011
R10077 dvss.t281 dvss.n744 76.1011
R10078 dvss.n1676 dvss.t584 76.1011
R10079 dvss.t335 dvss.n853 76.1011
R10080 dvss.t4 dvss.n3728 76.0887
R10081 dvss.t363 dvss.n3663 76.0887
R10082 dvss.t325 dvss.n2207 76.0887
R10083 dvss.t56 dvss.n2182 76.0887
R10084 dvss.t441 dvss.n2155 76.0887
R10085 dvss.t313 dvss.n2005 76.0887
R10086 dvss.t644 dvss.n1606 76.0887
R10087 dvss.t347 dvss.n1530 76.0887
R10088 dvss.n1183 dvss.t153 76.0887
R10089 dvss.n2258 dvss.t178 74.7229
R10090 dvss.t661 dvss.n3922 74.7229
R10091 dvss.t369 dvss.t169 74.6236
R10092 dvss.t169 dvss.t698 74.6236
R10093 dvss.t698 dvss.t526 74.6236
R10094 dvss.t526 dvss.t159 74.6236
R10095 dvss.t523 dvss.t382 74.6236
R10096 dvss.t168 dvss.t489 74.6236
R10097 dvss.t468 dvss.t168 74.6236
R10098 dvss.n4035 dvss.n4034 73.1255
R10099 dvss.n4034 dvss.n4033 73.1255
R10100 dvss.n4011 dvss.n3992 73.1255
R10101 dvss.n4012 dvss.n4011 73.1255
R10102 dvss.n3712 dvss 73.0358
R10103 dvss.n3774 dvss 73.0358
R10104 dvss.n3657 dvss 73.0358
R10105 dvss.n3672 dvss 73.0358
R10106 dvss.n2116 dvss 73.0358
R10107 dvss.n3017 dvss 73.0358
R10108 dvss.n2085 dvss 73.0358
R10109 dvss.n3067 dvss 73.0358
R10110 dvss.n2054 dvss 73.0358
R10111 dvss.n3117 dvss 73.0358
R10112 dvss.n1999 dvss 73.0358
R10113 dvss.n2014 dvss 73.0358
R10114 dvss.n1579 dvss 73.0358
R10115 dvss.n1639 dvss 73.0358
R10116 dvss.n1524 dvss 73.0358
R10117 dvss.n1539 dvss 73.0358
R10118 dvss.n1132 dvss 73.0358
R10119 dvss.n1140 dvss 73.0358
R10120 dvss dvss.n3857 73.0358
R10121 dvss.n3847 dvss 73.0358
R10122 dvss dvss.n3601 73.0358
R10123 dvss.n3591 dvss 73.0358
R10124 dvss dvss.n549 73.0358
R10125 dvss dvss.n3454 73.0358
R10126 dvss.n3333 dvss 73.0358
R10127 dvss dvss.n3335 73.0358
R10128 dvss dvss.n672 73.0358
R10129 dvss dvss.n3222 73.0358
R10130 dvss dvss.n1943 73.0358
R10131 dvss.n1933 dvss 73.0358
R10132 dvss dvss.n781 73.0358
R10133 dvss dvss.n1744 73.0358
R10134 dvss dvss.n1468 73.0358
R10135 dvss.n1458 dvss 73.0358
R10136 dvss dvss.n890 73.0358
R10137 dvss dvss.n1269 73.0358
R10138 dvss.n3990 dvss.n3989 66.9177
R10139 dvss.n3997 dvss.n3996 66.9014
R10140 dvss.n3999 dvss.n3995 66.9014
R10141 dvss.n4001 dvss.n3994 66.9014
R10142 dvss.n46 dvss.n45 66.771
R10143 dvss.n52 dvss.n47 66.771
R10144 dvss.n4003 dvss.n4002 66.6759
R10145 dvss.n429 dvss.t331 64.6673
R10146 dvss.n3562 dvss.t170 64.6673
R10147 dvss.n563 dvss.t534 64.6673
R10148 dvss.n3292 dvss.t196 64.6673
R10149 dvss.n687 dvss.t596 64.6673
R10150 dvss.n1862 dvss.t357 64.6673
R10151 dvss.n796 dvss.t559 64.6673
R10152 dvss.n1387 dvss.t561 64.6673
R10153 dvss.t355 dvss.n905 63.9189
R10154 dvss.n3902 dvss.t180 63.2272
R10155 dvss.t663 dvss.n328 63.2272
R10156 dvss.n329 dvss.n308 62.9701
R10157 dvss.n3809 dvss.n3808 62.9701
R10158 dvss.n3627 dvss.n3625 62.9701
R10159 dvss.n2199 dvss.n2198 62.9701
R10160 dvss.n2174 dvss.n2173 62.9701
R10161 dvss.n3152 dvss.n3151 62.9701
R10162 dvss.n1969 dvss.n1967 62.9701
R10163 dvss.n1674 dvss.n1673 62.9701
R10164 dvss.n1494 dvss.n1492 62.9701
R10165 dvss.n2889 dvss.t0 60.8054
R10166 dvss.t481 dvss.n4010 57.4543
R10167 dvss.n335 dvss.n334 57.0829
R10168 dvss.n3958 dvss.n337 57.0829
R10169 dvss.n386 dvss.n385 57.0829
R10170 dvss.n3882 dvss.n3880 57.0829
R10171 dvss.n520 dvss.n519 57.0829
R10172 dvss.n3507 dvss.n522 57.0829
R10173 dvss.n583 dvss.n582 57.0829
R10174 dvss.n3393 dvss.n585 57.0829
R10175 dvss.n646 dvss.n645 57.0829
R10176 dvss.n3276 dvss.n648 57.0829
R10177 dvss.n1841 dvss.n1840 57.0829
R10178 dvss.n1919 dvss.n1917 57.0829
R10179 dvss.n755 dvss.n754 57.0829
R10180 dvss.n1797 dvss.n757 57.0829
R10181 dvss.n1366 dvss.n1365 57.0829
R10182 dvss.n1444 dvss.n1442 57.0829
R10183 dvss.n864 dvss.n863 57.0829
R10184 dvss.n1322 dvss.n866 57.0829
R10185 dvss.n4083 dvss.n4082 57.0829
R10186 dvss.n4075 dvss.n4074 57.0829
R10187 dvss.n4117 dvss.n4115 57.0829
R10188 dvss.n270 dvss.n269 57.0829
R10189 dvss.n2981 dvss.n2288 57.0829
R10190 dvss.n2215 dvss.n2214 57.0829
R10191 dvss.n2309 dvss.n2308 57.0829
R10192 dvss.n2924 dvss.n2311 57.0829
R10193 dvss.n2645 dvss.n2644 57.0829
R10194 dvss.n2637 dvss.n2636 57.0829
R10195 dvss.n2692 dvss.n2691 57.0829
R10196 dvss.n2684 dvss.n2683 57.0829
R10197 dvss.n2739 dvss.n2738 57.0829
R10198 dvss.n2731 dvss.n2730 57.0829
R10199 dvss.n2786 dvss.n2785 57.0829
R10200 dvss.n2778 dvss.n2777 57.0829
R10201 dvss.n2833 dvss.n2832 57.0829
R10202 dvss.n2825 dvss.n2824 57.0829
R10203 dvss.n2257 dvss.t554 57.076
R10204 dvss.n2948 dvss.t696 57.076
R10205 dvss.t489 dvss.n4013 54.2898
R10206 dvss.n4014 dvss.t468 51.9608
R10207 dvss.t256 dvss.n2237 49.9195
R10208 dvss.n2916 dvss.t113 49.9195
R10209 dvss.n3941 dvss.t214 48.4282
R10210 dvss.t133 dvss.n456 48.4282
R10211 dvss.t28 dvss.n3496 48.4282
R10212 dvss.n3384 dvss.t42 48.4282
R10213 dvss.t295 dvss.n3264 48.4282
R10214 dvss.t569 dvss.n1909 48.4282
R10215 dvss.t279 dvss.n1786 48.4282
R10216 dvss.t586 dvss.n1434 48.4282
R10217 dvss.t337 dvss.n1311 48.4282
R10218 dvss.n4032 dvss.t369 47.3803
R10219 dvss.n3792 dvss.n3706 46.2505
R10220 dvss.n3783 dvss.n3713 46.2505
R10221 dvss.n495 dvss.n494 46.2505
R10222 dvss.n486 dvss.n485 46.2505
R10223 dvss.n3035 dvss.n2111 46.2505
R10224 dvss.n3026 dvss.n2117 46.2505
R10225 dvss.n3085 dvss.n2080 46.2505
R10226 dvss.n3076 dvss.n2086 46.2505
R10227 dvss.n3135 dvss.n2048 46.2505
R10228 dvss.n3126 dvss.n2055 46.2505
R10229 dvss.n731 dvss.n730 46.2505
R10230 dvss.n722 dvss.n721 46.2505
R10231 dvss.n1657 dvss.n1573 46.2505
R10232 dvss.n1648 dvss.n1580 46.2505
R10233 dvss.n840 dvss.n839 46.2505
R10234 dvss.n831 dvss.n830 46.2505
R10235 dvss.n1129 dvss.n1128 46.2505
R10236 dvss.n1137 dvss.n1136 46.2505
R10237 dvss.n412 dvss.n411 46.2505
R10238 dvss.n414 dvss.n413 46.2505
R10239 dvss.n3533 dvss.n3532 46.2505
R10240 dvss.n3535 dvss.n3534 46.2505
R10241 dvss.n3436 dvss.n3432 46.2505
R10242 dvss.n3453 dvss.n3452 46.2505
R10243 dvss.n617 dvss.n616 46.2505
R10244 dvss.n3339 dvss.n3334 46.2505
R10245 dvss.n3207 dvss.n3206 46.2505
R10246 dvss.n3221 dvss.n3220 46.2505
R10247 dvss.n1823 dvss.n1822 46.2505
R10248 dvss.n1825 dvss.n1824 46.2505
R10249 dvss.n1729 dvss.n1728 46.2505
R10250 dvss.n1743 dvss.n1742 46.2505
R10251 dvss.n1348 dvss.n1347 46.2505
R10252 dvss.n1350 dvss.n1349 46.2505
R10253 dvss.n1254 dvss.n1253 46.2505
R10254 dvss.n1268 dvss.n1267 46.2505
R10255 dvss.n237 dvss.n236 45.0005
R10256 dvss.n57 dvss.n43 45.0005
R10257 dvss.t307 dvss.n43 45.0005
R10258 dvss.n44 dvss.n42 45.0005
R10259 dvss.t307 dvss.n42 45.0005
R10260 dvss.n134 dvss.n133 45.0005
R10261 dvss.n174 dvss.n173 45.0005
R10262 dvss.n3774 dvss 44.424
R10263 dvss.n3672 dvss 44.424
R10264 dvss.n3017 dvss 44.424
R10265 dvss.n3067 dvss 44.424
R10266 dvss.n3117 dvss 44.424
R10267 dvss.n2014 dvss 44.424
R10268 dvss.n1639 dvss 44.424
R10269 dvss.n1539 dvss 44.424
R10270 dvss.n1140 dvss 44.424
R10271 dvss.n3847 dvss 44.424
R10272 dvss.n3591 dvss 44.424
R10273 dvss.n3454 dvss 44.424
R10274 dvss.n3335 dvss 44.424
R10275 dvss.n3222 dvss 44.424
R10276 dvss.n1933 dvss 44.424
R10277 dvss.n1744 dvss 44.424
R10278 dvss.n1458 dvss 44.424
R10279 dvss.n1269 dvss 44.424
R10280 dvss.t237 dvss.n1022 43.2419
R10281 dvss.t249 dvss.n2413 43.2419
R10282 dvss.n2987 dvss.t260 39.2225
R10283 dvss.t109 dvss.n600 39.2225
R10284 dvss.n3931 dvss.t208 38.0508
R10285 dvss.n3896 dvss.t127 38.0508
R10286 dvss.n2987 dvss.t32 38.0508
R10287 dvss.t38 dvss.n600 38.0508
R10288 dvss.n2158 dvss.t301 38.0508
R10289 dvss.n1898 dvss.t573 38.0508
R10290 dvss.n1609 dvss.t289 38.0508
R10291 dvss.n1423 dvss.t592 38.0508
R10292 dvss.n1124 dvss.t343 38.0508
R10293 dvss.n1098 dvss.t232 37.7206
R10294 dvss.n1020 dvss.t253 37.7206
R10295 dvss.t159 dvss.n4031 37.3121
R10296 dvss.n4031 dvss.t382 37.3121
R10297 dvss.n234 dvss.n233 36.563
R10298 dvss.t501 dvss.t374 36.1649
R10299 dvss.n1229 dvss.n1228 36.1417
R10300 dvss.n1228 dvss.n1227 36.1417
R10301 dvss.n1227 dvss.n1061 36.1417
R10302 dvss.n1221 dvss.n1061 36.1417
R10303 dvss.n1221 dvss.n1220 36.1417
R10304 dvss.n1220 dvss.n1219 36.1417
R10305 dvss.n1219 dvss.n1069 36.1417
R10306 dvss.n1212 dvss.n1069 36.1417
R10307 dvss.n1212 dvss.n1211 36.1417
R10308 dvss.n1211 dvss.n1210 36.1417
R10309 dvss.n1210 dvss.n1080 36.1417
R10310 dvss.n1204 dvss.n1080 36.1417
R10311 dvss.n1204 dvss.n1203 36.1417
R10312 dvss.n1203 dvss.n1202 36.1417
R10313 dvss.n1202 dvss.n1093 36.1417
R10314 dvss.n1196 dvss.n1093 36.1417
R10315 dvss.n1195 dvss.n1194 36.1417
R10316 dvss.n1194 dvss.n1106 36.1417
R10317 dvss.n1188 dvss.n1106 36.1417
R10318 dvss.n1188 dvss.n1187 36.1417
R10319 dvss.n1187 dvss.n1186 36.1417
R10320 dvss.n1186 dvss.n1113 36.1417
R10321 dvss.n1180 dvss.n1113 36.1417
R10322 dvss.n1180 dvss.n1179 36.1417
R10323 dvss.n1179 dvss.n1178 36.1417
R10324 dvss.n1178 dvss.n1120 36.1417
R10325 dvss.n1172 dvss.n1120 36.1417
R10326 dvss.n1172 dvss.n1171 36.1417
R10327 dvss.n1171 dvss.n1170 36.1417
R10328 dvss.n1170 dvss.n1148 36.1417
R10329 dvss.n1164 dvss.n1148 36.1417
R10330 dvss.n1164 dvss.n1163 36.1417
R10331 dvss.n1163 dvss.n850 36.1417
R10332 dvss.n1496 dvss.n850 36.1417
R10333 dvss.n1496 dvss.n849 36.1417
R10334 dvss.n1501 dvss.n849 36.1417
R10335 dvss.n1501 dvss.n846 36.1417
R10336 dvss.n1507 dvss.n846 36.1417
R10337 dvss.n1507 dvss.n845 36.1417
R10338 dvss.n1513 dvss.n845 36.1417
R10339 dvss.n1513 dvss.n841 36.1417
R10340 dvss.n1519 dvss.n841 36.1417
R10341 dvss.n1519 dvss.n837 36.1417
R10342 dvss.n1528 dvss.n837 36.1417
R10343 dvss.n1528 dvss.n833 36.1417
R10344 dvss.n1535 dvss.n833 36.1417
R10345 dvss.n1535 dvss.n827 36.1417
R10346 dvss.n1543 dvss.n827 36.1417
R10347 dvss.n1543 dvss.n824 36.1417
R10348 dvss.n1550 dvss.n824 36.1417
R10349 dvss.n1550 dvss.n819 36.1417
R10350 dvss.n1558 dvss.n819 36.1417
R10351 dvss.n1558 dvss.n816 36.1417
R10352 dvss.n1564 dvss.n816 36.1417
R10353 dvss.n1564 dvss.n814 36.1417
R10354 dvss.n1671 dvss.n814 36.1417
R10355 dvss.n1671 dvss.n815 36.1417
R10356 dvss.n1667 dvss.n815 36.1417
R10357 dvss.n1667 dvss.n1666 36.1417
R10358 dvss.n1666 dvss.n1569 36.1417
R10359 dvss.n1662 dvss.n1569 36.1417
R10360 dvss.n1662 dvss.n1661 36.1417
R10361 dvss.n1661 dvss.n1572 36.1417
R10362 dvss.n1575 dvss.n1572 36.1417
R10363 dvss.n1653 dvss.n1575 36.1417
R10364 dvss.n1653 dvss.n1652 36.1417
R10365 dvss.n1652 dvss.n1578 36.1417
R10366 dvss.n1644 dvss.n1578 36.1417
R10367 dvss.n1644 dvss.n1643 36.1417
R10368 dvss.n1643 dvss.n1584 36.1417
R10369 dvss.n1636 dvss.n1584 36.1417
R10370 dvss.n1636 dvss.n1635 36.1417
R10371 dvss.n1635 dvss.n1588 36.1417
R10372 dvss.n1592 dvss.n1588 36.1417
R10373 dvss.n1626 dvss.n1592 36.1417
R10374 dvss.n1626 dvss.n1625 36.1417
R10375 dvss.n1625 dvss.n741 36.1417
R10376 dvss.n1971 dvss.n741 36.1417
R10377 dvss.n1971 dvss.n740 36.1417
R10378 dvss.n1976 dvss.n740 36.1417
R10379 dvss.n1976 dvss.n737 36.1417
R10380 dvss.n1982 dvss.n737 36.1417
R10381 dvss.n1982 dvss.n736 36.1417
R10382 dvss.n1988 dvss.n736 36.1417
R10383 dvss.n1988 dvss.n732 36.1417
R10384 dvss.n1994 dvss.n732 36.1417
R10385 dvss.n1994 dvss.n728 36.1417
R10386 dvss.n2003 dvss.n728 36.1417
R10387 dvss.n2003 dvss.n724 36.1417
R10388 dvss.n2010 dvss.n724 36.1417
R10389 dvss.n2010 dvss.n718 36.1417
R10390 dvss.n2018 dvss.n718 36.1417
R10391 dvss.n2018 dvss.n715 36.1417
R10392 dvss.n2025 dvss.n715 36.1417
R10393 dvss.n2025 dvss.n710 36.1417
R10394 dvss.n2033 dvss.n710 36.1417
R10395 dvss.n2033 dvss.n707 36.1417
R10396 dvss.n2039 dvss.n707 36.1417
R10397 dvss.n2039 dvss.n705 36.1417
R10398 dvss.n3149 dvss.n705 36.1417
R10399 dvss.n3149 dvss.n706 36.1417
R10400 dvss.n3145 dvss.n706 36.1417
R10401 dvss.n3145 dvss.n3144 36.1417
R10402 dvss.n3144 dvss.n2044 36.1417
R10403 dvss.n3140 dvss.n2044 36.1417
R10404 dvss.n3140 dvss.n3139 36.1417
R10405 dvss.n3139 dvss.n2047 36.1417
R10406 dvss.n2050 dvss.n2047 36.1417
R10407 dvss.n3131 dvss.n2050 36.1417
R10408 dvss.n3131 dvss.n3130 36.1417
R10409 dvss.n3130 dvss.n2053 36.1417
R10410 dvss.n3122 dvss.n2053 36.1417
R10411 dvss.n3122 dvss.n3121 36.1417
R10412 dvss.n3121 dvss.n2059 36.1417
R10413 dvss.n3114 dvss.n2059 36.1417
R10414 dvss.n3114 dvss.n3113 36.1417
R10415 dvss.n3113 dvss.n2063 36.1417
R10416 dvss.n2067 dvss.n2063 36.1417
R10417 dvss.n3104 dvss.n2067 36.1417
R10418 dvss.n3104 dvss.n3103 36.1417
R10419 dvss.n3103 dvss.n2070 36.1417
R10420 dvss.n3099 dvss.n2070 36.1417
R10421 dvss.n3099 dvss.n3098 36.1417
R10422 dvss.n3098 dvss.n2073 36.1417
R10423 dvss.n3094 dvss.n2073 36.1417
R10424 dvss.n3094 dvss.n3093 36.1417
R10425 dvss.n3093 dvss.n2076 36.1417
R10426 dvss.n3089 dvss.n2076 36.1417
R10427 dvss.n3089 dvss.n3088 36.1417
R10428 dvss.n3088 dvss.n2079 36.1417
R10429 dvss.n3081 dvss.n2079 36.1417
R10430 dvss.n3081 dvss.n3080 36.1417
R10431 dvss.n3080 dvss.n2084 36.1417
R10432 dvss.n3072 dvss.n2084 36.1417
R10433 dvss.n3072 dvss.n3071 36.1417
R10434 dvss.n3071 dvss.n2090 36.1417
R10435 dvss.n3064 dvss.n2090 36.1417
R10436 dvss.n3064 dvss.n3063 36.1417
R10437 dvss.n3063 dvss.n2094 36.1417
R10438 dvss.n2098 dvss.n2094 36.1417
R10439 dvss.n3054 dvss.n2098 36.1417
R10440 dvss.n3054 dvss.n3053 36.1417
R10441 dvss.n3053 dvss.n2101 36.1417
R10442 dvss.n3049 dvss.n2101 36.1417
R10443 dvss.n3049 dvss.n3048 36.1417
R10444 dvss.n3048 dvss.n2104 36.1417
R10445 dvss.n3044 dvss.n2104 36.1417
R10446 dvss.n3044 dvss.n3043 36.1417
R10447 dvss.n3043 dvss.n2107 36.1417
R10448 dvss.n3039 dvss.n2107 36.1417
R10449 dvss.n3039 dvss.n3038 36.1417
R10450 dvss.n3038 dvss.n2110 36.1417
R10451 dvss.n3031 dvss.n2110 36.1417
R10452 dvss.n3031 dvss.n3030 36.1417
R10453 dvss.n3030 dvss.n2115 36.1417
R10454 dvss.n3022 dvss.n2115 36.1417
R10455 dvss.n3022 dvss.n3021 36.1417
R10456 dvss.n3021 dvss.n2121 36.1417
R10457 dvss.n3014 dvss.n2121 36.1417
R10458 dvss.n3014 dvss.n3013 36.1417
R10459 dvss.n3013 dvss.n2125 36.1417
R10460 dvss.n2129 dvss.n2125 36.1417
R10461 dvss.n3004 dvss.n2129 36.1417
R10462 dvss.n3004 dvss.n3003 36.1417
R10463 dvss.n3003 dvss.n505 36.1417
R10464 dvss.n3629 dvss.n505 36.1417
R10465 dvss.n3629 dvss.n504 36.1417
R10466 dvss.n3634 dvss.n504 36.1417
R10467 dvss.n3634 dvss.n501 36.1417
R10468 dvss.n3640 dvss.n501 36.1417
R10469 dvss.n3640 dvss.n500 36.1417
R10470 dvss.n3646 dvss.n500 36.1417
R10471 dvss.n3646 dvss.n496 36.1417
R10472 dvss.n3652 dvss.n496 36.1417
R10473 dvss.n3652 dvss.n492 36.1417
R10474 dvss.n3661 dvss.n492 36.1417
R10475 dvss.n3661 dvss.n488 36.1417
R10476 dvss.n3668 dvss.n488 36.1417
R10477 dvss.n3668 dvss.n482 36.1417
R10478 dvss.n3676 dvss.n482 36.1417
R10479 dvss.n3676 dvss.n479 36.1417
R10480 dvss.n3683 dvss.n479 36.1417
R10481 dvss.n3683 dvss.n474 36.1417
R10482 dvss.n3691 dvss.n474 36.1417
R10483 dvss.n3691 dvss.n471 36.1417
R10484 dvss.n3697 dvss.n471 36.1417
R10485 dvss.n3697 dvss.n469 36.1417
R10486 dvss.n3806 dvss.n469 36.1417
R10487 dvss.n3806 dvss.n470 36.1417
R10488 dvss.n3802 dvss.n470 36.1417
R10489 dvss.n3802 dvss.n3801 36.1417
R10490 dvss.n3801 dvss.n3702 36.1417
R10491 dvss.n3797 dvss.n3702 36.1417
R10492 dvss.n3797 dvss.n3796 36.1417
R10493 dvss.n3796 dvss.n3705 36.1417
R10494 dvss.n3708 dvss.n3705 36.1417
R10495 dvss.n3788 dvss.n3708 36.1417
R10496 dvss.n3788 dvss.n3787 36.1417
R10497 dvss.n3787 dvss.n3711 36.1417
R10498 dvss.n3779 dvss.n3711 36.1417
R10499 dvss.n3779 dvss.n3778 36.1417
R10500 dvss.n3778 dvss.n3733 36.1417
R10501 dvss.n3771 dvss.n3733 36.1417
R10502 dvss.n3771 dvss.n3770 36.1417
R10503 dvss.n3770 dvss.n3737 36.1417
R10504 dvss.n3741 dvss.n3737 36.1417
R10505 dvss.n3761 dvss.n3741 36.1417
R10506 dvss.n3761 dvss.n3760 36.1417
R10507 dvss.n3760 dvss.n3756 36.1417
R10508 dvss.n3756 dvss.n311 36.1417
R10509 dvss.n4051 dvss.n311 36.1417
R10510 dvss.n4051 dvss.n312 36.1417
R10511 dvss.n4047 dvss.n312 36.1417
R10512 dvss.n963 dvss.n962 36.1417
R10513 dvss.n962 dvss.n960 36.1417
R10514 dvss.n969 dvss.n960 36.1417
R10515 dvss.n973 dvss.n969 36.1417
R10516 dvss.n975 dvss.n973 36.1417
R10517 dvss.n975 dvss.n957 36.1417
R10518 dvss.n981 dvss.n957 36.1417
R10519 dvss.n988 dvss.n981 36.1417
R10520 dvss.n990 dvss.n988 36.1417
R10521 dvss.n990 dvss.n954 36.1417
R10522 dvss.n996 dvss.n954 36.1417
R10523 dvss.n1010 dvss.n996 36.1417
R10524 dvss.n1012 dvss.n1010 36.1417
R10525 dvss.n1012 dvss.n935 36.1417
R10526 dvss.n1017 dvss.n935 36.1417
R10527 dvss.n1017 dvss.n936 36.1417
R10528 dvss.n949 dvss.n936 36.1417
R10529 dvss.n949 dvss.n902 36.1417
R10530 dvss.n902 dvss.n900 36.1417
R10531 dvss.n1245 dvss.n900 36.1417
R10532 dvss.n1245 dvss.n896 36.1417
R10533 dvss.n1258 dvss.n896 36.1417
R10534 dvss.n1258 dvss.n888 36.1417
R10535 dvss.n1273 dvss.n888 36.1417
R10536 dvss.n1274 dvss.n1273 36.1417
R10537 dvss.n1274 dvss.n885 36.1417
R10538 dvss.n885 dvss.n879 36.1417
R10539 dvss.n1294 dvss.n879 36.1417
R10540 dvss.n1295 dvss.n1294 36.1417
R10541 dvss.n1295 dvss.n875 36.1417
R10542 dvss.n875 dvss.n867 36.1417
R10543 dvss.n872 dvss.n867 36.1417
R10544 dvss.n1315 dvss.n872 36.1417
R10545 dvss.n1315 dvss.n858 36.1417
R10546 dvss.n1488 dvss.n858 36.1417
R10547 dvss.n1488 dvss.n859 36.1417
R10548 dvss.n1330 dvss.n859 36.1417
R10549 dvss.n1331 dvss.n1330 36.1417
R10550 dvss.n1335 dvss.n1331 36.1417
R10551 dvss.n1336 dvss.n1335 36.1417
R10552 dvss.n1401 dvss.n1336 36.1417
R10553 dvss.n1401 dvss.n1340 36.1417
R10554 dvss.n1345 dvss.n1340 36.1417
R10555 dvss.n1408 dvss.n1345 36.1417
R10556 dvss.n1411 dvss.n1408 36.1417
R10557 dvss.n1411 dvss.n1351 36.1417
R10558 dvss.n1356 dvss.n1351 36.1417
R10559 dvss.n1357 dvss.n1356 36.1417
R10560 dvss.n1378 dvss.n1357 36.1417
R10561 dvss.n1378 dvss.n1360 36.1417
R10562 dvss.n1368 dvss.n1360 36.1417
R10563 dvss.n1369 dvss.n1368 36.1417
R10564 dvss.n1377 dvss.n1369 36.1417
R10565 dvss.n1377 dvss.n1373 36.1417
R10566 dvss.n1373 dvss.n807 36.1417
R10567 dvss.n1678 dvss.n807 36.1417
R10568 dvss.n1678 dvss.n802 36.1417
R10569 dvss.n1705 dvss.n802 36.1417
R10570 dvss.n1705 dvss.n803 36.1417
R10571 dvss.n1692 dvss.n803 36.1417
R10572 dvss.n1698 dvss.n1692 36.1417
R10573 dvss.n1698 dvss.n793 36.1417
R10574 dvss.n793 dvss.n791 36.1417
R10575 dvss.n1720 dvss.n791 36.1417
R10576 dvss.n1720 dvss.n787 36.1417
R10577 dvss.n1733 dvss.n787 36.1417
R10578 dvss.n1733 dvss.n779 36.1417
R10579 dvss.n1748 dvss.n779 36.1417
R10580 dvss.n1749 dvss.n1748 36.1417
R10581 dvss.n1749 dvss.n776 36.1417
R10582 dvss.n776 dvss.n770 36.1417
R10583 dvss.n1769 dvss.n770 36.1417
R10584 dvss.n1770 dvss.n1769 36.1417
R10585 dvss.n1770 dvss.n766 36.1417
R10586 dvss.n766 dvss.n758 36.1417
R10587 dvss.n763 dvss.n758 36.1417
R10588 dvss.n1790 dvss.n763 36.1417
R10589 dvss.n1790 dvss.n749 36.1417
R10590 dvss.n1963 dvss.n749 36.1417
R10591 dvss.n1963 dvss.n750 36.1417
R10592 dvss.n1805 dvss.n750 36.1417
R10593 dvss.n1806 dvss.n1805 36.1417
R10594 dvss.n1810 dvss.n1806 36.1417
R10595 dvss.n1811 dvss.n1810 36.1417
R10596 dvss.n1876 dvss.n1811 36.1417
R10597 dvss.n1876 dvss.n1815 36.1417
R10598 dvss.n1820 dvss.n1815 36.1417
R10599 dvss.n1883 dvss.n1820 36.1417
R10600 dvss.n1886 dvss.n1883 36.1417
R10601 dvss.n1886 dvss.n1826 36.1417
R10602 dvss.n1831 dvss.n1826 36.1417
R10603 dvss.n1832 dvss.n1831 36.1417
R10604 dvss.n1853 dvss.n1832 36.1417
R10605 dvss.n1853 dvss.n1835 36.1417
R10606 dvss.n1843 dvss.n1835 36.1417
R10607 dvss.n1844 dvss.n1843 36.1417
R10608 dvss.n1852 dvss.n1844 36.1417
R10609 dvss.n1852 dvss.n1848 36.1417
R10610 dvss.n1848 dvss.n698 36.1417
R10611 dvss.n3156 dvss.n698 36.1417
R10612 dvss.n3156 dvss.n693 36.1417
R10613 dvss.n3183 dvss.n693 36.1417
R10614 dvss.n3183 dvss.n694 36.1417
R10615 dvss.n3170 dvss.n694 36.1417
R10616 dvss.n3176 dvss.n3170 36.1417
R10617 dvss.n3176 dvss.n684 36.1417
R10618 dvss.n684 dvss.n682 36.1417
R10619 dvss.n3198 dvss.n682 36.1417
R10620 dvss.n3198 dvss.n678 36.1417
R10621 dvss.n3211 dvss.n678 36.1417
R10622 dvss.n3211 dvss.n670 36.1417
R10623 dvss.n3226 dvss.n670 36.1417
R10624 dvss.n3227 dvss.n3226 36.1417
R10625 dvss.n3227 dvss.n667 36.1417
R10626 dvss.n667 dvss.n661 36.1417
R10627 dvss.n3247 dvss.n661 36.1417
R10628 dvss.n3248 dvss.n3247 36.1417
R10629 dvss.n3248 dvss.n657 36.1417
R10630 dvss.n657 dvss.n649 36.1417
R10631 dvss.n654 dvss.n649 36.1417
R10632 dvss.n3269 dvss.n654 36.1417
R10633 dvss.n3269 dvss.n640 36.1417
R10634 dvss.n3284 dvss.n640 36.1417
R10635 dvss.n3284 dvss.n634 36.1417
R10636 dvss.n3303 dvss.n634 36.1417
R10637 dvss.n3303 dvss.n635 36.1417
R10638 dvss.n635 dvss.n628 36.1417
R10639 dvss.n3309 dvss.n628 36.1417
R10640 dvss.n3309 dvss.n623 36.1417
R10641 dvss.n3320 dvss.n623 36.1417
R10642 dvss.n3320 dvss.n618 36.1417
R10643 dvss.n3329 dvss.n618 36.1417
R10644 dvss.n3329 dvss.n613 36.1417
R10645 dvss.n3346 dvss.n613 36.1417
R10646 dvss.n3346 dvss.n606 36.1417
R10647 dvss.n3353 dvss.n606 36.1417
R10648 dvss.n3353 dvss.n602 36.1417
R10649 dvss.n3363 dvss.n602 36.1417
R10650 dvss.n3363 dvss.n597 36.1417
R10651 dvss.n3377 dvss.n597 36.1417
R10652 dvss.n3377 dvss.n586 36.1417
R10653 dvss.n3386 dvss.n586 36.1417
R10654 dvss.n3386 dvss.n580 36.1417
R10655 dvss.n3398 dvss.n580 36.1417
R10656 dvss.n3399 dvss.n3398 36.1417
R10657 dvss.n3399 dvss.n575 36.1417
R10658 dvss.n575 dvss.n568 36.1417
R10659 dvss.n569 dvss.n568 36.1417
R10660 dvss.n3412 dvss.n569 36.1417
R10661 dvss.n3412 dvss.n559 36.1417
R10662 dvss.n3430 dvss.n559 36.1417
R10663 dvss.n3431 dvss.n3430 36.1417
R10664 dvss.n3431 dvss.n556 36.1417
R10665 dvss.n556 dvss.n550 36.1417
R10666 dvss.n550 dvss.n545 36.1417
R10667 dvss.n3462 dvss.n545 36.1417
R10668 dvss.n3462 dvss.n546 36.1417
R10669 dvss.n546 dvss.n541 36.1417
R10670 dvss.n541 dvss.n535 36.1417
R10671 dvss.n3479 dvss.n535 36.1417
R10672 dvss.n3480 dvss.n3479 36.1417
R10673 dvss.n3480 dvss.n531 36.1417
R10674 dvss.n531 dvss.n523 36.1417
R10675 dvss.n528 dvss.n523 36.1417
R10676 dvss.n3500 dvss.n528 36.1417
R10677 dvss.n3500 dvss.n514 36.1417
R10678 dvss.n3621 dvss.n514 36.1417
R10679 dvss.n3621 dvss.n515 36.1417
R10680 dvss.n3515 dvss.n515 36.1417
R10681 dvss.n3516 dvss.n3515 36.1417
R10682 dvss.n3520 dvss.n3516 36.1417
R10683 dvss.n3521 dvss.n3520 36.1417
R10684 dvss.n3552 dvss.n3521 36.1417
R10685 dvss.n3552 dvss.n3525 36.1417
R10686 dvss.n3530 dvss.n3525 36.1417
R10687 dvss.n3548 dvss.n3530 36.1417
R10688 dvss.n3551 dvss.n3548 36.1417
R10689 dvss.n3551 dvss.n3536 36.1417
R10690 dvss.n3541 dvss.n3536 36.1417
R10691 dvss.n3585 dvss.n3541 36.1417
R10692 dvss.n3585 dvss.n374 36.1417
R10693 dvss.n3893 dvss.n374 36.1417
R10694 dvss.n3893 dvss.n375 36.1417
R10695 dvss.n379 dvss.n375 36.1417
R10696 dvss.n452 dvss.n379 36.1417
R10697 dvss.n454 dvss.n452 36.1417
R10698 dvss.n454 dvss.n441 36.1417
R10699 dvss.n462 dvss.n441 36.1417
R10700 dvss.n462 dvss.n388 36.1417
R10701 dvss.n393 dvss.n388 36.1417
R10702 dvss.n394 dvss.n393 36.1417
R10703 dvss.n395 dvss.n394 36.1417
R10704 dvss.n399 dvss.n395 36.1417
R10705 dvss.n400 dvss.n399 36.1417
R10706 dvss.n3819 dvss.n400 36.1417
R10707 dvss.n3819 dvss.n404 36.1417
R10708 dvss.n409 dvss.n404 36.1417
R10709 dvss.n3826 dvss.n409 36.1417
R10710 dvss.n3829 dvss.n3826 36.1417
R10711 dvss.n3829 dvss.n415 36.1417
R10712 dvss.n420 dvss.n415 36.1417
R10713 dvss.n421 dvss.n420 36.1417
R10714 dvss.n421 dvss.n348 36.1417
R10715 dvss.n3934 dvss.n348 36.1417
R10716 dvss.n3934 dvss.n342 36.1417
R10717 dvss.n3945 dvss.n342 36.1417
R10718 dvss.n3945 dvss.n338 36.1417
R10719 dvss.n338 dvss.n333 36.1417
R10720 dvss.n3964 dvss.n333 36.1417
R10721 dvss.n3964 dvss.n323 36.1417
R10722 dvss.n3973 dvss.n323 36.1417
R10723 dvss.n3973 dvss.n319 36.1417
R10724 dvss.n3979 dvss.n319 36.1417
R10725 dvss.n3979 dvss.n313 36.1417
R10726 dvss.n1055 dvss.n1054 36.1417
R10727 dvss.n1054 dvss.n1053 36.1417
R10728 dvss.n1053 dvss.n917 36.1417
R10729 dvss.n1048 dvss.n917 36.1417
R10730 dvss.n1048 dvss.n1047 36.1417
R10731 dvss.n1047 dvss.n1046 36.1417
R10732 dvss.n1046 dvss.n922 36.1417
R10733 dvss.n1040 dvss.n922 36.1417
R10734 dvss.n1040 dvss.n1039 36.1417
R10735 dvss.n1039 dvss.n1038 36.1417
R10736 dvss.n1038 dvss.n927 36.1417
R10737 dvss.n1032 dvss.n927 36.1417
R10738 dvss.n1032 dvss.n1031 36.1417
R10739 dvss.n1031 dvss.n1030 36.1417
R10740 dvss.n1030 dvss.n932 36.1417
R10741 dvss.n946 dvss.n932 36.1417
R10742 dvss.n1237 dvss.n903 36.1417
R10743 dvss.n1237 dvss.n1236 36.1417
R10744 dvss.n1236 dvss.n897 36.1417
R10745 dvss.n1250 dvss.n897 36.1417
R10746 dvss.n1250 dvss.n891 36.1417
R10747 dvss.n1263 dvss.n891 36.1417
R10748 dvss.n1263 dvss.n887 36.1417
R10749 dvss.n1277 dvss.n887 36.1417
R10750 dvss.n1277 dvss.n882 36.1417
R10751 dvss.n1287 dvss.n882 36.1417
R10752 dvss.n1287 dvss.n878 36.1417
R10753 dvss.n1304 dvss.n878 36.1417
R10754 dvss.n1304 dvss.n869 36.1417
R10755 dvss.n1319 dvss.n869 36.1417
R10756 dvss.n1319 dvss.n1318 36.1417
R10757 dvss.n1318 dvss.n861 36.1417
R10758 dvss.n1327 dvss.n861 36.1417
R10759 dvss.n1486 dvss.n1327 36.1417
R10760 dvss.n1486 dvss.n1485 36.1417
R10761 dvss.n1485 dvss.n1329 36.1417
R10762 dvss.n1481 dvss.n1329 36.1417
R10763 dvss.n1480 dvss.n1334 36.1417
R10764 dvss.n1341 dvss.n1334 36.1417
R10765 dvss.n1473 dvss.n1341 36.1417
R10766 dvss.n1473 dvss.n1472 36.1417
R10767 dvss.n1472 dvss.n1344 36.1417
R10768 dvss.n1352 dvss.n1344 36.1417
R10769 dvss.n1464 dvss.n1352 36.1417
R10770 dvss.n1464 dvss.n1463 36.1417
R10771 dvss.n1463 dvss.n1355 36.1417
R10772 dvss.n1361 dvss.n1355 36.1417
R10773 dvss.n1453 dvss.n1361 36.1417
R10774 dvss.n1453 dvss.n1452 36.1417
R10775 dvss.n1452 dvss.n1364 36.1417
R10776 dvss.n1374 dvss.n1364 36.1417
R10777 dvss.n1439 dvss.n1374 36.1417
R10778 dvss.n1439 dvss.n1438 36.1417
R10779 dvss.n1438 dvss.n804 36.1417
R10780 dvss.n1684 dvss.n804 36.1417
R10781 dvss.n1703 dvss.n1684 36.1417
R10782 dvss.n1703 dvss.n1702 36.1417
R10783 dvss.n1702 dvss.n1691 36.1417
R10784 dvss.n1712 dvss.n794 36.1417
R10785 dvss.n1712 dvss.n1711 36.1417
R10786 dvss.n1711 dvss.n788 36.1417
R10787 dvss.n1725 dvss.n788 36.1417
R10788 dvss.n1725 dvss.n782 36.1417
R10789 dvss.n1738 dvss.n782 36.1417
R10790 dvss.n1738 dvss.n778 36.1417
R10791 dvss.n1752 dvss.n778 36.1417
R10792 dvss.n1752 dvss.n773 36.1417
R10793 dvss.n1762 dvss.n773 36.1417
R10794 dvss.n1762 dvss.n769 36.1417
R10795 dvss.n1779 dvss.n769 36.1417
R10796 dvss.n1779 dvss.n760 36.1417
R10797 dvss.n1794 dvss.n760 36.1417
R10798 dvss.n1794 dvss.n1793 36.1417
R10799 dvss.n1793 dvss.n752 36.1417
R10800 dvss.n1802 dvss.n752 36.1417
R10801 dvss.n1961 dvss.n1802 36.1417
R10802 dvss.n1961 dvss.n1960 36.1417
R10803 dvss.n1960 dvss.n1804 36.1417
R10804 dvss.n1956 dvss.n1804 36.1417
R10805 dvss.n1955 dvss.n1809 36.1417
R10806 dvss.n1816 dvss.n1809 36.1417
R10807 dvss.n1948 dvss.n1816 36.1417
R10808 dvss.n1948 dvss.n1947 36.1417
R10809 dvss.n1947 dvss.n1819 36.1417
R10810 dvss.n1827 dvss.n1819 36.1417
R10811 dvss.n1939 dvss.n1827 36.1417
R10812 dvss.n1939 dvss.n1938 36.1417
R10813 dvss.n1938 dvss.n1830 36.1417
R10814 dvss.n1836 dvss.n1830 36.1417
R10815 dvss.n1928 dvss.n1836 36.1417
R10816 dvss.n1928 dvss.n1927 36.1417
R10817 dvss.n1927 dvss.n1839 36.1417
R10818 dvss.n1849 dvss.n1839 36.1417
R10819 dvss.n1914 dvss.n1849 36.1417
R10820 dvss.n1914 dvss.n1913 36.1417
R10821 dvss.n1913 dvss.n695 36.1417
R10822 dvss.n3162 dvss.n695 36.1417
R10823 dvss.n3181 dvss.n3162 36.1417
R10824 dvss.n3181 dvss.n3180 36.1417
R10825 dvss.n3180 dvss.n3169 36.1417
R10826 dvss.n3190 dvss.n685 36.1417
R10827 dvss.n3190 dvss.n3189 36.1417
R10828 dvss.n3189 dvss.n679 36.1417
R10829 dvss.n3203 dvss.n679 36.1417
R10830 dvss.n3203 dvss.n673 36.1417
R10831 dvss.n3216 dvss.n673 36.1417
R10832 dvss.n3216 dvss.n669 36.1417
R10833 dvss.n3230 dvss.n669 36.1417
R10834 dvss.n3230 dvss.n664 36.1417
R10835 dvss.n3240 dvss.n664 36.1417
R10836 dvss.n3240 dvss.n660 36.1417
R10837 dvss.n3257 dvss.n660 36.1417
R10838 dvss.n3257 dvss.n651 36.1417
R10839 dvss.n3273 dvss.n651 36.1417
R10840 dvss.n3273 dvss.n3272 36.1417
R10841 dvss.n3272 dvss.n643 36.1417
R10842 dvss.n3281 dvss.n643 36.1417
R10843 dvss.n3282 dvss.n3281 36.1417
R10844 dvss.n3282 dvss.n636 36.1417
R10845 dvss.n3301 dvss.n636 36.1417
R10846 dvss.n3301 dvss.n3300 36.1417
R10847 dvss.n3297 dvss.n626 36.1417
R10848 dvss.n3317 dvss.n626 36.1417
R10849 dvss.n3318 dvss.n3317 36.1417
R10850 dvss.n3318 dvss.n621 36.1417
R10851 dvss.n621 dvss.n614 36.1417
R10852 dvss.n3343 dvss.n614 36.1417
R10853 dvss.n3344 dvss.n3343 36.1417
R10854 dvss.n3344 dvss.n604 36.1417
R10855 dvss.n3355 dvss.n604 36.1417
R10856 dvss.n3356 dvss.n3355 36.1417
R10857 dvss.n3356 dvss.n598 36.1417
R10858 dvss.n3368 dvss.n598 36.1417
R10859 dvss.n3368 dvss.n588 36.1417
R10860 dvss.n3390 dvss.n588 36.1417
R10861 dvss.n3390 dvss.n3389 36.1417
R10862 dvss.n3389 dvss.n591 36.1417
R10863 dvss.n591 dvss.n578 36.1417
R10864 dvss.n3402 dvss.n578 36.1417
R10865 dvss.n3402 dvss.n566 36.1417
R10866 dvss.n3416 dvss.n566 36.1417
R10867 dvss.n3416 dvss.n567 36.1417
R10868 dvss.n3422 dvss.n561 36.1417
R10869 dvss.n3422 dvss.n558 36.1417
R10870 dvss.n3439 dvss.n558 36.1417
R10871 dvss.n3439 dvss.n551 36.1417
R10872 dvss.n3447 dvss.n551 36.1417
R10873 dvss.n3447 dvss.n547 36.1417
R10874 dvss.n3460 dvss.n547 36.1417
R10875 dvss.n3460 dvss.n3459 36.1417
R10876 dvss.n3459 dvss.n538 36.1417
R10877 dvss.n3472 dvss.n538 36.1417
R10878 dvss.n3472 dvss.n534 36.1417
R10879 dvss.n3489 dvss.n534 36.1417
R10880 dvss.n3489 dvss.n525 36.1417
R10881 dvss.n3504 dvss.n525 36.1417
R10882 dvss.n3504 dvss.n3503 36.1417
R10883 dvss.n3503 dvss.n517 36.1417
R10884 dvss.n3512 dvss.n517 36.1417
R10885 dvss.n3619 dvss.n3512 36.1417
R10886 dvss.n3619 dvss.n3618 36.1417
R10887 dvss.n3618 dvss.n3514 36.1417
R10888 dvss.n3614 dvss.n3514 36.1417
R10889 dvss.n3613 dvss.n3519 36.1417
R10890 dvss.n3526 dvss.n3519 36.1417
R10891 dvss.n3606 dvss.n3526 36.1417
R10892 dvss.n3606 dvss.n3605 36.1417
R10893 dvss.n3605 dvss.n3529 36.1417
R10894 dvss.n3537 dvss.n3529 36.1417
R10895 dvss.n3597 dvss.n3537 36.1417
R10896 dvss.n3597 dvss.n3596 36.1417
R10897 dvss.n3596 dvss.n3540 36.1417
R10898 dvss.n3540 dvss.n376 36.1417
R10899 dvss.n3891 dvss.n376 36.1417
R10900 dvss.n3891 dvss.n3890 36.1417
R10901 dvss.n3890 dvss.n378 36.1417
R10902 dvss.n448 dvss.n378 36.1417
R10903 dvss.n448 dvss.n442 36.1417
R10904 dvss.n459 dvss.n442 36.1417
R10905 dvss.n459 dvss.n389 36.1417
R10906 dvss.n3875 dvss.n389 36.1417
R10907 dvss.n3875 dvss.n3874 36.1417
R10908 dvss.n3874 dvss.n392 36.1417
R10909 dvss.n3870 dvss.n392 36.1417
R10910 dvss.n3869 dvss.n398 36.1417
R10911 dvss.n405 dvss.n398 36.1417
R10912 dvss.n3862 dvss.n405 36.1417
R10913 dvss.n3862 dvss.n3861 36.1417
R10914 dvss.n3861 dvss.n408 36.1417
R10915 dvss.n416 dvss.n408 36.1417
R10916 dvss.n3853 dvss.n416 36.1417
R10917 dvss.n3853 dvss.n3852 36.1417
R10918 dvss.n3852 dvss.n419 36.1417
R10919 dvss.n3841 dvss.n419 36.1417
R10920 dvss.n3841 dvss.n347 36.1417
R10921 dvss.n3938 dvss.n347 36.1417
R10922 dvss.n3938 dvss.n340 36.1417
R10923 dvss.n3955 dvss.n340 36.1417
R10924 dvss.n3955 dvss.n3954 36.1417
R10925 dvss.n3954 dvss.n331 36.1417
R10926 dvss.n331 dvss.n320 36.1417
R10927 dvss.n3975 dvss.n320 36.1417
R10928 dvss.n3976 dvss.n3975 36.1417
R10929 dvss.n3976 dvss.n314 36.1417
R10930 dvss.n3984 dvss.n314 36.1417
R10931 dvss.n2887 dvss.n2392 36.1417
R10932 dvss.n2884 dvss.n2392 36.1417
R10933 dvss.n2884 dvss.n2883 36.1417
R10934 dvss.n2883 dvss.n2395 36.1417
R10935 dvss.n2879 dvss.n2395 36.1417
R10936 dvss.n2879 dvss.n2878 36.1417
R10937 dvss.n2878 dvss.n2400 36.1417
R10938 dvss.n2874 dvss.n2400 36.1417
R10939 dvss.n2874 dvss.n2873 36.1417
R10940 dvss.n2873 dvss.n2403 36.1417
R10941 dvss.n2866 dvss.n2403 36.1417
R10942 dvss.n2866 dvss.n2865 36.1417
R10943 dvss.n2865 dvss.n2411 36.1417
R10944 dvss.n2416 dvss.n2411 36.1417
R10945 dvss.n2858 dvss.n2416 36.1417
R10946 dvss.n2858 dvss.n2857 36.1417
R10947 dvss.n2854 dvss.n2853 36.1417
R10948 dvss.n2853 dvss.n2423 36.1417
R10949 dvss.n2847 dvss.n2423 36.1417
R10950 dvss.n2847 dvss.n2846 36.1417
R10951 dvss.n2846 dvss.n2429 36.1417
R10952 dvss.n2842 dvss.n2429 36.1417
R10953 dvss.n2842 dvss.n2841 36.1417
R10954 dvss.n2841 dvss.n2434 36.1417
R10955 dvss.n2837 dvss.n2434 36.1417
R10956 dvss.n2837 dvss.n2836 36.1417
R10957 dvss.n2836 dvss.n2437 36.1417
R10958 dvss.n2829 dvss.n2437 36.1417
R10959 dvss.n2829 dvss.n2828 36.1417
R10960 dvss.n2828 dvss.n2444 36.1417
R10961 dvss.n2821 dvss.n2444 36.1417
R10962 dvss.n2821 dvss.n2820 36.1417
R10963 dvss.n2820 dvss.n2448 36.1417
R10964 dvss.n2813 dvss.n2448 36.1417
R10965 dvss.n2813 dvss.n2812 36.1417
R10966 dvss.n2812 dvss.n2453 36.1417
R10967 dvss.n2808 dvss.n2453 36.1417
R10968 dvss.n2807 dvss.n2456 36.1417
R10969 dvss.n2462 dvss.n2456 36.1417
R10970 dvss.n2800 dvss.n2462 36.1417
R10971 dvss.n2800 dvss.n2799 36.1417
R10972 dvss.n2799 dvss.n2465 36.1417
R10973 dvss.n2795 dvss.n2465 36.1417
R10974 dvss.n2795 dvss.n2794 36.1417
R10975 dvss.n2794 dvss.n2470 36.1417
R10976 dvss.n2790 dvss.n2470 36.1417
R10977 dvss.n2790 dvss.n2789 36.1417
R10978 dvss.n2789 dvss.n2473 36.1417
R10979 dvss.n2782 dvss.n2473 36.1417
R10980 dvss.n2782 dvss.n2781 36.1417
R10981 dvss.n2781 dvss.n2480 36.1417
R10982 dvss.n2774 dvss.n2480 36.1417
R10983 dvss.n2774 dvss.n2773 36.1417
R10984 dvss.n2773 dvss.n2484 36.1417
R10985 dvss.n2766 dvss.n2484 36.1417
R10986 dvss.n2766 dvss.n2765 36.1417
R10987 dvss.n2765 dvss.n2489 36.1417
R10988 dvss.n2761 dvss.n2489 36.1417
R10989 dvss.n2760 dvss.n2492 36.1417
R10990 dvss.n2498 dvss.n2492 36.1417
R10991 dvss.n2753 dvss.n2498 36.1417
R10992 dvss.n2753 dvss.n2752 36.1417
R10993 dvss.n2752 dvss.n2501 36.1417
R10994 dvss.n2748 dvss.n2501 36.1417
R10995 dvss.n2748 dvss.n2747 36.1417
R10996 dvss.n2747 dvss.n2506 36.1417
R10997 dvss.n2743 dvss.n2506 36.1417
R10998 dvss.n2743 dvss.n2742 36.1417
R10999 dvss.n2742 dvss.n2509 36.1417
R11000 dvss.n2735 dvss.n2509 36.1417
R11001 dvss.n2735 dvss.n2734 36.1417
R11002 dvss.n2734 dvss.n2516 36.1417
R11003 dvss.n2727 dvss.n2516 36.1417
R11004 dvss.n2727 dvss.n2726 36.1417
R11005 dvss.n2726 dvss.n2520 36.1417
R11006 dvss.n2719 dvss.n2520 36.1417
R11007 dvss.n2719 dvss.n2718 36.1417
R11008 dvss.n2718 dvss.n2525 36.1417
R11009 dvss.n2714 dvss.n2525 36.1417
R11010 dvss.n2713 dvss.n2528 36.1417
R11011 dvss.n2534 dvss.n2528 36.1417
R11012 dvss.n2706 dvss.n2534 36.1417
R11013 dvss.n2706 dvss.n2705 36.1417
R11014 dvss.n2705 dvss.n2537 36.1417
R11015 dvss.n2701 dvss.n2537 36.1417
R11016 dvss.n2701 dvss.n2700 36.1417
R11017 dvss.n2700 dvss.n2542 36.1417
R11018 dvss.n2696 dvss.n2542 36.1417
R11019 dvss.n2696 dvss.n2695 36.1417
R11020 dvss.n2695 dvss.n2545 36.1417
R11021 dvss.n2688 dvss.n2545 36.1417
R11022 dvss.n2688 dvss.n2687 36.1417
R11023 dvss.n2687 dvss.n2552 36.1417
R11024 dvss.n2680 dvss.n2552 36.1417
R11025 dvss.n2680 dvss.n2679 36.1417
R11026 dvss.n2679 dvss.n2556 36.1417
R11027 dvss.n2672 dvss.n2556 36.1417
R11028 dvss.n2672 dvss.n2671 36.1417
R11029 dvss.n2671 dvss.n2561 36.1417
R11030 dvss.n2667 dvss.n2561 36.1417
R11031 dvss.n2666 dvss.n2564 36.1417
R11032 dvss.n2570 dvss.n2564 36.1417
R11033 dvss.n2659 dvss.n2570 36.1417
R11034 dvss.n2659 dvss.n2658 36.1417
R11035 dvss.n2658 dvss.n2573 36.1417
R11036 dvss.n2654 dvss.n2573 36.1417
R11037 dvss.n2654 dvss.n2653 36.1417
R11038 dvss.n2653 dvss.n2578 36.1417
R11039 dvss.n2649 dvss.n2578 36.1417
R11040 dvss.n2649 dvss.n2648 36.1417
R11041 dvss.n2648 dvss.n2581 36.1417
R11042 dvss.n2641 dvss.n2581 36.1417
R11043 dvss.n2641 dvss.n2640 36.1417
R11044 dvss.n2640 dvss.n2588 36.1417
R11045 dvss.n2633 dvss.n2588 36.1417
R11046 dvss.n2633 dvss.n2632 36.1417
R11047 dvss.n2632 dvss.n2592 36.1417
R11048 dvss.n2625 dvss.n2592 36.1417
R11049 dvss.n2625 dvss.n2624 36.1417
R11050 dvss.n2624 dvss.n2597 36.1417
R11051 dvss.n2620 dvss.n2597 36.1417
R11052 dvss.n2619 dvss.n2600 36.1417
R11053 dvss.n2606 dvss.n2600 36.1417
R11054 dvss.n2612 dvss.n2606 36.1417
R11055 dvss.n2612 dvss.n2611 36.1417
R11056 dvss.n2611 dvss.n2323 36.1417
R11057 dvss.n2892 dvss.n2323 36.1417
R11058 dvss.n2892 dvss.n2322 36.1417
R11059 dvss.n2897 dvss.n2322 36.1417
R11060 dvss.n2897 dvss.n2318 36.1417
R11061 dvss.n2903 dvss.n2318 36.1417
R11062 dvss.n2903 dvss.n2317 36.1417
R11063 dvss.n2910 dvss.n2317 36.1417
R11064 dvss.n2910 dvss.n2312 36.1417
R11065 dvss.n2921 dvss.n2312 36.1417
R11066 dvss.n2921 dvss.n2920 36.1417
R11067 dvss.n2920 dvss.n2307 36.1417
R11068 dvss.n2931 dvss.n2307 36.1417
R11069 dvss.n2931 dvss.n2304 36.1417
R11070 dvss.n2938 dvss.n2304 36.1417
R11071 dvss.n2938 dvss.n2303 36.1417
R11072 dvss.n2943 dvss.n2303 36.1417
R11073 dvss.n2950 dvss.n2299 36.1417
R11074 dvss.n2950 dvss.n2297 36.1417
R11075 dvss.n2959 dvss.n2297 36.1417
R11076 dvss.n2959 dvss.n2294 36.1417
R11077 dvss.n2965 dvss.n2294 36.1417
R11078 dvss.n2965 dvss.n2293 36.1417
R11079 dvss.n2970 dvss.n2293 36.1417
R11080 dvss.n2970 dvss.n2289 36.1417
R11081 dvss.n2977 dvss.n2289 36.1417
R11082 dvss.n2977 dvss.n2212 36.1417
R11083 dvss.n2984 dvss.n2212 36.1417
R11084 dvss.n2984 dvss.n2213 36.1417
R11085 dvss.n2227 dvss.n2213 36.1417
R11086 dvss.n2227 dvss.n2221 36.1417
R11087 dvss.n2235 dvss.n2221 36.1417
R11088 dvss.n2235 dvss.n2222 36.1417
R11089 dvss.n2222 dvss.n2217 36.1417
R11090 dvss.n2283 dvss.n2217 36.1417
R11091 dvss.n2283 dvss.n2282 36.1417
R11092 dvss.n2282 dvss.n2243 36.1417
R11093 dvss.n2278 dvss.n2243 36.1417
R11094 dvss.n2277 dvss.n2246 36.1417
R11095 dvss.n2270 dvss.n2246 36.1417
R11096 dvss.n2270 dvss.n259 36.1417
R11097 dvss.n4131 dvss.n259 36.1417
R11098 dvss.n4131 dvss.n4130 36.1417
R11099 dvss.n4130 dvss.n262 36.1417
R11100 dvss.n4126 dvss.n262 36.1417
R11101 dvss.n4126 dvss.n4125 36.1417
R11102 dvss.n4125 dvss.n265 36.1417
R11103 dvss.n4121 dvss.n265 36.1417
R11104 dvss.n4121 dvss.n4120 36.1417
R11105 dvss.n4120 dvss.n268 36.1417
R11106 dvss.n367 dvss.n268 36.1417
R11107 dvss.n367 dvss.n357 36.1417
R11108 dvss.n361 dvss.n357 36.1417
R11109 dvss.n361 dvss.n351 36.1417
R11110 dvss.n351 dvss.n272 36.1417
R11111 dvss.n4110 dvss.n272 36.1417
R11112 dvss.n4110 dvss.n4109 36.1417
R11113 dvss.n4109 dvss.n275 36.1417
R11114 dvss.n4105 dvss.n275 36.1417
R11115 dvss.n4104 dvss.n278 36.1417
R11116 dvss.n282 dvss.n278 36.1417
R11117 dvss.n4097 dvss.n282 36.1417
R11118 dvss.n4097 dvss.n4096 36.1417
R11119 dvss.n4096 dvss.n285 36.1417
R11120 dvss.n4092 dvss.n285 36.1417
R11121 dvss.n4092 dvss.n4091 36.1417
R11122 dvss.n4091 dvss.n288 36.1417
R11123 dvss.n4087 dvss.n288 36.1417
R11124 dvss.n4087 dvss.n4086 36.1417
R11125 dvss.n4086 dvss.n291 36.1417
R11126 dvss.n4079 dvss.n291 36.1417
R11127 dvss.n4079 dvss.n4078 36.1417
R11128 dvss.n4078 dvss.n296 36.1417
R11129 dvss.n4071 dvss.n296 36.1417
R11130 dvss.n4071 dvss.n4070 36.1417
R11131 dvss.n4070 dvss.n300 36.1417
R11132 dvss.n4063 dvss.n300 36.1417
R11133 dvss.n4063 dvss.n4062 36.1417
R11134 dvss.n4062 dvss.n303 36.1417
R11135 dvss.n4058 dvss.n303 36.1417
R11136 dvss.n1196 dvss.n1195 35.7652
R11137 dvss.n2224 dvss.t254 35.6569
R11138 dvss.t111 dvss.n2314 35.6569
R11139 dvss.t212 dvss.n345 34.5917
R11140 dvss.n445 dvss.t123 34.5917
R11141 dvss.t26 dvss.n532 34.5917
R11142 dvss.t40 dvss.n594 34.5917
R11143 dvss.t299 dvss.n658 34.5917
R11144 dvss.n1902 dvss.t565 34.5917
R11145 dvss.t287 dvss.n767 34.5917
R11146 dvss.n1427 dvss.t590 34.5917
R11147 dvss.t341 dvss.n876 34.5917
R11148 dvss.n3766 dvss 33.9483
R11149 dvss.n3687 dvss 33.9483
R11150 dvss.n3009 dvss 33.9483
R11151 dvss.n3059 dvss 33.9483
R11152 dvss.n3109 dvss 33.9483
R11153 dvss.n2029 dvss 33.9483
R11154 dvss.n1631 dvss 33.9483
R11155 dvss.n1554 dvss 33.9483
R11156 dvss.n1157 dvss 33.9483
R11157 dvss.n3950 dvss 33.9483
R11158 dvss.n3886 dvss 33.9483
R11159 dvss.n3485 dvss 33.9483
R11160 dvss.n3374 dvss 33.9483
R11161 dvss.n3253 dvss 33.9483
R11162 dvss.n1923 dvss 33.9483
R11163 dvss.n1775 dvss 33.9483
R11164 dvss.n1448 dvss 33.9483
R11165 dvss.n1300 dvss 33.9483
R11166 dvss.n3925 dvss.t667 32.1345
R11167 dvss.t184 dvss.n3898 32.1345
R11168 dvss.n3909 dvss.t227 31.6138
R11169 dvss.t206 dvss.t669 31.1326
R11170 dvss.t131 dvss.t176 31.1326
R11171 dvss.t34 dvss.t258 31.1326
R11172 dvss.t115 dvss.t46 31.1326
R11173 dvss.t297 dvss.t539 31.1326
R11174 dvss.t571 dvss.t575 31.1326
R11175 dvss.t285 dvss.t529 31.1326
R11176 dvss.t588 dvss.t198 31.1326
R11177 dvss.t339 dvss.t239 31.1326
R11178 dvss.n1085 dvss.n1084 30.6481
R11179 dvss.n999 dvss.n998 30.6481
R11180 dvss.t174 dvss.n370 28.7399
R11181 dvss.t665 dvss.n3930 28.7399
R11182 dvss.n401 dvss.t429 28.1205
R11183 dvss.n3522 dvss.t537 28.1205
R11184 dvss.n3425 dvss.t436 28.1205
R11185 dvss.n3312 dvss.t595 28.1205
R11186 dvss.n3193 dvss.t173 28.1205
R11187 dvss.n1812 dvss.t122 28.1205
R11188 dvss.n1715 dvss.t733 28.1205
R11189 dvss.n1337 dvss.t15 28.1205
R11190 dvss.n1240 dvss.t13 28.1205
R11191 dvss.n279 dvss.t230 28.1205
R11192 dvss.n2247 dvss.t557 28.1205
R11193 dvss.n2953 dvss.t467 28.1205
R11194 dvss.n2601 dvss.t731 28.1205
R11195 dvss.n2565 dvss.t381 28.1205
R11196 dvss.n2529 dvss.t224 28.1205
R11197 dvss.n2493 dvss.t545 28.1205
R11198 dvss.n2457 dvss.t494 28.1205
R11199 dvss.n2424 dvss.t100 28.1205
R11200 dvss.n3837 dvss.n422 27.2737
R11201 dvss.n3583 dvss.n3582 27.2737
R11202 dvss.n3467 dvss.n3466 27.2737
R11203 dvss.n3351 dvss.n3350 27.2737
R11204 dvss.n3235 dvss.n3234 27.2737
R11205 dvss.n1894 dvss.n1855 27.2737
R11206 dvss.n1757 dvss.n1756 27.2737
R11207 dvss.n1419 dvss.n1380 27.2737
R11208 dvss.n1282 dvss.n1281 27.2737
R11209 dvss.n911 dvss.t200 26.6829
R11210 dvss.n3 dvss.t104 24.9236
R11211 dvss.n3 dvss.t108 24.9236
R11212 dvss.n218 dvss.t551 24.9236
R11213 dvss.n218 dvss.t549 24.9236
R11214 dvss.n99 dvss.t165 24.9236
R11215 dvss.n99 dvss.t161 24.9236
R11216 dvss.n113 dvss.t720 24.9236
R11217 dvss.n113 dvss.t710 24.9236
R11218 dvss.n115 dvss.t722 24.9236
R11219 dvss.n115 dvss.t702 24.9236
R11220 dvss.n110 dvss.t726 24.9236
R11221 dvss.n110 dvss.t728 24.9236
R11222 dvss.n124 dvss.t716 24.9236
R11223 dvss.n124 dvss.t706 24.9236
R11224 dvss.n107 dvss.t712 24.9236
R11225 dvss.n107 dvss.t730 24.9236
R11226 dvss.n104 dvss.t714 24.9236
R11227 dvss.n104 dvss.t700 24.9236
R11228 dvss.n103 dvss.t724 24.9236
R11229 dvss.n103 dvss.t704 24.9236
R11230 dvss.n7 dvss.t306 24.9236
R11231 dvss.n7 dvss.t518 24.9236
R11232 dvss.n21 dvss.t71 24.9236
R11233 dvss.n21 dvss.t93 24.9236
R11234 dvss.n23 dvss.t73 24.9236
R11235 dvss.n23 dvss.t85 24.9236
R11236 dvss.n18 dvss.t77 24.9236
R11237 dvss.n18 dvss.t79 24.9236
R11238 dvss.n32 dvss.t67 24.9236
R11239 dvss.n32 dvss.t89 24.9236
R11240 dvss.n15 dvss.t63 24.9236
R11241 dvss.n15 dvss.t81 24.9236
R11242 dvss.n12 dvss.t65 24.9236
R11243 dvss.n12 dvss.t83 24.9236
R11244 dvss.n11 dvss.t75 24.9236
R11245 dvss.n11 dvss.t87 24.9236
R11246 dvss.n96 dvss.t452 24.9236
R11247 dvss.n96 dvss.t448 24.9236
R11248 dvss.n70 dvss.t391 24.9236
R11249 dvss.n70 dvss.t413 24.9236
R11250 dvss.n69 dvss.t393 24.9236
R11251 dvss.n69 dvss.t405 24.9236
R11252 dvss.n77 dvss.t397 24.9236
R11253 dvss.n77 dvss.t399 24.9236
R11254 dvss.n66 dvss.t387 24.9236
R11255 dvss.n66 dvss.t409 24.9236
R11256 dvss.n86 dvss.t415 24.9236
R11257 dvss.n86 dvss.t401 24.9236
R11258 dvss.n63 dvss.t417 24.9236
R11259 dvss.n63 dvss.t403 24.9236
R11260 dvss.n92 dvss.t395 24.9236
R11261 dvss.n92 dvss.t407 24.9236
R11262 dvss.n190 dvss.t603 24.9236
R11263 dvss.n190 dvss.t627 24.9236
R11264 dvss.n192 dvss.t617 24.9236
R11265 dvss.n192 dvss.t629 24.9236
R11266 dvss.n187 dvss.t609 24.9236
R11267 dvss.n187 dvss.t623 24.9236
R11268 dvss.n201 dvss.t613 24.9236
R11269 dvss.n201 dvss.t599 24.9236
R11270 dvss.n184 dvss.t615 24.9236
R11271 dvss.n184 dvss.t601 24.9236
R11272 dvss.n210 dvss.t605 24.9236
R11273 dvss.n210 dvss.t619 24.9236
R11274 dvss.n181 dvss.t607 24.9236
R11275 dvss.n181 dvss.t621 24.9236
R11276 dvss.n1005 dvss.n1003 22.5639
R11277 dvss.n2406 dvss.n2404 22.5639
R11278 dvss.t135 dvss.n3822 22.5415
R11279 dvss.n3570 dvss.t469 22.5415
R11280 dvss.t186 dvss.n3441 22.5415
R11281 dvss.t16 dvss.n3322 22.5415
R11282 dvss.t636 dvss.n3200 22.5415
R11283 dvss.t462 dvss.n1879 22.5415
R11284 dvss.t679 dvss.n1722 22.5415
R11285 dvss.t511 dvss.n1404 22.5415
R11286 dvss.t426 dvss.n1247 22.5415
R11287 dvss.n4045 dvss.n4039 22.2727
R11288 dvss.n1098 dvss.t278 22.0013
R11289 dvss.n1020 dvss.t375 22.0013
R11290 dvss.n3767 dvss.n3766 21.8222
R11291 dvss.n3687 dvss.n3686 21.8222
R11292 dvss.n3010 dvss.n3009 21.8222
R11293 dvss.n3060 dvss.n3059 21.8222
R11294 dvss.n3110 dvss.n3109 21.8222
R11295 dvss.n2029 dvss.n2028 21.8222
R11296 dvss.n1632 dvss.n1631 21.8222
R11297 dvss.n1554 dvss.n1553 21.8222
R11298 dvss.n1157 dvss.n1152 21.8222
R11299 dvss.n3950 dvss.n3947 21.8222
R11300 dvss.n3887 dvss.n3886 21.8222
R11301 dvss.n3486 dvss.n3485 21.8222
R11302 dvss.n3375 dvss.n3374 21.8222
R11303 dvss.n3254 dvss.n3253 21.8222
R11304 dvss.n1924 dvss.n1923 21.8222
R11305 dvss.n1776 dvss.n1775 21.8222
R11306 dvss.n1449 dvss.n1448 21.8222
R11307 dvss.n1301 dvss.n1300 21.8222
R11308 dvss.n401 dvss.t332 21.2805
R11309 dvss.n3522 dvss.t171 21.2805
R11310 dvss.n3425 dvss.t535 21.2805
R11311 dvss.n3312 dvss.t197 21.2805
R11312 dvss.n3193 dvss.t597 21.2805
R11313 dvss.n1812 dvss.t358 21.2805
R11314 dvss.n1715 dvss.t560 21.2805
R11315 dvss.n1337 dvss.t562 21.2805
R11316 dvss.n1240 dvss.t356 21.2805
R11317 dvss.n1004 dvss.t238 21.2805
R11318 dvss.n1004 dvss.t236 21.2805
R11319 dvss.n279 dvss.t228 21.2805
R11320 dvss.n2247 dvss.t555 21.2805
R11321 dvss.n2953 dvss.t697 21.2805
R11322 dvss.n2601 dvss.t270 21.2805
R11323 dvss.n2565 dvss.t434 21.2805
R11324 dvss.n2529 dvss.t1 21.2805
R11325 dvss.n2493 dvss.t558 21.2805
R11326 dvss.n2457 dvss.t455 21.2805
R11327 dvss.n2424 dvss.t658 21.2805
R11328 dvss.n2405 dvss.t251 21.2805
R11329 dvss.n2405 dvss.t250 21.2805
R11330 dvss.n1022 dvss.t99 20.3576
R11331 dvss.n2413 dvss.t267 20.3576
R11332 dvss.n4013 dvss.t523 20.3343
R11333 dvss.n3739 dvss.t217 20.0005
R11334 dvss.n3739 dvss.t51 20.0005
R11335 dvss.n475 dvss.t126 20.0005
R11336 dvss.n475 dvss.t498 20.0005
R11337 dvss.n2127 dvss.t31 20.0005
R11338 dvss.n2127 dvss.t226 20.0005
R11339 dvss.n2096 dvss.t45 20.0005
R11340 dvss.n2096 dvss.t310 20.0005
R11341 dvss.n2065 dvss.t294 20.0005
R11342 dvss.n2065 dvss.t525 20.0005
R11343 dvss.n711 dvss.t564 20.0005
R11344 dvss.n711 dvss.t493 20.0005
R11345 dvss.n1590 dvss.t284 20.0005
R11346 dvss.n1590 dvss.t431 20.0005
R11347 dvss.n820 dvss.t583 20.0005
R11348 dvss.n820 dvss.t522 20.0005
R11349 dvss.n1153 dvss.t334 20.0005
R11350 dvss.n1153 dvss.t373 20.0005
R11351 dvss.n3948 dvss.t670 20.0005
R11352 dvss.n3948 dvss.t500 20.0005
R11353 dvss.n381 dvss.t177 20.0005
R11354 dvss.n381 dvss.t496 20.0005
R11355 dvss.n3483 dvss.t259 20.0005
R11356 dvss.n3483 dvss.t520 20.0005
R11357 dvss.n3372 dvss.t116 20.0005
R11358 dvss.n3372 dvss.t371 20.0005
R11359 dvss.n3251 dvss.t540 20.0005
R11360 dvss.n3251 dvss.t97 20.0005
R11361 dvss.n1846 dvss.t576 20.0005
R11362 dvss.n1846 dvss.t641 20.0005
R11363 dvss.n1773 dvss.t530 20.0005
R11364 dvss.n1773 dvss.t514 20.0005
R11365 dvss.n1371 dvss.t199 20.0005
R11366 dvss.n1371 dvss.t433 20.0005
R11367 dvss.n1298 dvss.t240 20.0005
R11368 dvss.n1298 dvss.t491 20.0005
R11369 dvss.n429 dvss.n428 18.8324
R11370 dvss.n3562 dvss.n3561 18.8324
R11371 dvss.n573 dvss.n563 18.8324
R11372 dvss.n3292 dvss.n631 18.8324
R11373 dvss.n3186 dvss.n687 18.8324
R11374 dvss.n1862 dvss.n1861 18.8324
R11375 dvss.n1708 dvss.n796 18.8324
R11376 dvss.n1387 dvss.n1386 18.8324
R11377 dvss.n1199 dvss.t231 18.6559
R11378 dvss.n1233 dvss.n905 18.6144
R11379 dvss.n3730 dvss.t6 18.3666
R11380 dvss.n3666 dvss.t365 18.3666
R11381 dvss.n2988 dvss.t327 18.3666
R11382 dvss.n2184 dvss.t58 18.3666
R11383 dvss.n2159 dvss.t439 18.3666
R11384 dvss.n2008 dvss.t319 18.3666
R11385 dvss.n1610 dvss.t642 18.3666
R11386 dvss.n1533 dvss.t353 18.3666
R11387 dvss.n1122 dvss.t157 18.3666
R11388 dvss.n946 dvss 18.0711
R11389 dvss.n1481 dvss 18.0711
R11390 dvss dvss.n1480 18.0711
R11391 dvss.n1691 dvss 18.0711
R11392 dvss dvss.n794 18.0711
R11393 dvss.n1956 dvss 18.0711
R11394 dvss dvss.n1955 18.0711
R11395 dvss.n3169 dvss 18.0711
R11396 dvss dvss.n685 18.0711
R11397 dvss.n3300 dvss 18.0711
R11398 dvss.n3297 dvss 18.0711
R11399 dvss.n567 dvss 18.0711
R11400 dvss dvss.n561 18.0711
R11401 dvss.n3614 dvss 18.0711
R11402 dvss dvss.n3613 18.0711
R11403 dvss.n3870 dvss 18.0711
R11404 dvss dvss.n3869 18.0711
R11405 dvss.n3984 dvss 18.0711
R11406 dvss.n2857 dvss 18.0711
R11407 dvss.n2854 dvss 18.0711
R11408 dvss.n2808 dvss 18.0711
R11409 dvss dvss.n2807 18.0711
R11410 dvss.n2761 dvss 18.0711
R11411 dvss dvss.n2760 18.0711
R11412 dvss.n2714 dvss 18.0711
R11413 dvss dvss.n2713 18.0711
R11414 dvss.n2667 dvss 18.0711
R11415 dvss dvss.n2666 18.0711
R11416 dvss.n2620 dvss 18.0711
R11417 dvss dvss.n2619 18.0711
R11418 dvss.n2943 dvss 18.0711
R11419 dvss dvss.n2299 18.0711
R11420 dvss.n2278 dvss 18.0711
R11421 dvss dvss.n2277 18.0711
R11422 dvss.n4105 dvss 18.0711
R11423 dvss dvss.n4104 18.0711
R11424 dvss.n4058 dvss 18.0711
R11425 dvss.n4002 dvss.t695 18.0005
R11426 dvss dvss.n903 17.6946
R11427 dvss.n3996 dvss.t146 17.4005
R11428 dvss.n3996 dvss.t683 17.4005
R11429 dvss.n3995 dvss.t657 17.4005
R11430 dvss.n3995 dvss.t686 17.4005
R11431 dvss.n3994 dvss.t148 17.4005
R11432 dvss.n3994 dvss.t482 17.4005
R11433 dvss.n4002 dvss.t487 17.4005
R11434 dvss.n3989 dvss.t689 17.4005
R11435 dvss.n3989 dvss.t385 17.4005
R11436 dvss.n45 dvss.t95 17.4005
R11437 dvss.n45 dvss.t692 17.4005
R11438 dvss.n47 dvss.t308 17.4005
R11439 dvss.n47 dvss.t221 17.4005
R11440 dvss.n3897 dvss.n352 17.2441
R11441 dvss.n121 dvss.n111 16.3561
R11442 dvss.n126 dvss.n123 16.3561
R11443 dvss.n130 dvss.n108 16.3561
R11444 dvss.n141 dvss.n140 16.3561
R11445 dvss.n146 dvss.n144 16.3561
R11446 dvss.n150 dvss.n100 16.3561
R11447 dvss.n151 dvss.n150 16.3561
R11448 dvss.n79 dvss.n76 16.3561
R11449 dvss.n83 dvss.n67 16.3561
R11450 dvss.n88 dvss.n85 16.3561
R11451 dvss.n167 dvss.n166 16.3561
R11452 dvss.n163 dvss.n162 16.3561
R11453 dvss.n159 dvss.n158 16.3561
R11454 dvss.n158 dvss.n157 16.3561
R11455 dvss.n4024 dvss.n4023 16.3427
R11456 dvss.n3834 dvss.n3833 16.2668
R11457 dvss.n3581 dvss.n3546 16.2668
R11458 dvss.n3465 dvss.n542 16.2668
R11459 dvss.n3349 dvss.n609 16.2668
R11460 dvss.n3233 dvss.n3232 16.2668
R11461 dvss.n1891 dvss.n1890 16.2668
R11462 dvss.n1755 dvss.n1754 16.2668
R11463 dvss.n1416 dvss.n1415 16.2668
R11464 dvss.n1280 dvss.n1279 16.2668
R11465 dvss.n4025 dvss.n4024 16.1789
R11466 dvss.n117 dvss.n114 16.1783
R11467 dvss.n74 dvss.n71 16.1783
R11468 dvss.n29 dvss.n19 16.132
R11469 dvss.n34 dvss.n31 16.132
R11470 dvss.n38 dvss.n16 16.132
R11471 dvss.n244 dvss.n243 16.132
R11472 dvss.n249 dvss.n247 16.132
R11473 dvss.n253 dvss.n8 16.132
R11474 dvss.n254 dvss.n253 16.132
R11475 dvss.n1214 dvss.t268 15.9908
R11476 dvss.n25 dvss.n22 15.9567
R11477 dvss.n139 dvss.n138 15.8227
R11478 dvss.n169 dvss.n168 15.8227
R11479 dvss.n2889 dvss.n2320 15.7029
R11480 dvss.n135 dvss.n134 15.6449
R11481 dvss.n173 dvss.n172 15.6449
R11482 dvss.n4021 dvss.n3987 15.6268
R11483 dvss.n242 dvss.n241 15.606
R11484 dvss.n152 dvss.n151 15.2894
R11485 dvss.n157 dvss.n97 15.2894
R11486 dvss.n911 dvss.t246 15.1155
R11487 dvss.n255 dvss.n254 15.08
R11488 dvss.n145 dvss.n100 14.9338
R11489 dvss.n159 dvss.n94 14.9338
R11490 dvss.n248 dvss.n8 14.7293
R11491 dvss.n198 dvss.n188 14.7205
R11492 dvss.n203 dvss.n200 14.7205
R11493 dvss.n207 dvss.n185 14.7205
R11494 dvss.n212 dvss.n209 14.7205
R11495 dvss.n231 dvss.n182 14.7205
R11496 dvss.n227 dvss.n226 14.7205
R11497 dvss.n223 dvss.n222 14.7205
R11498 dvss.n222 dvss.n221 14.7205
R11499 dvss.n4142 dvss.n2 14.7205
R11500 dvss.n4140 dvss.n4139 14.7205
R11501 dvss.n4139 dvss.n4 14.7205
R11502 dvss.n194 dvss.n191 14.5605
R11503 dvss.n238 dvss.n237 14.5539
R11504 dvss.n138 dvss.n105 14.0449
R11505 dvss.n141 dvss.n101 14.0449
R11506 dvss.n169 dvss.n64 14.0449
R11507 dvss.n166 dvss.n93 14.0449
R11508 dvss.n4022 dvss.n4021 13.9386
R11509 dvss.n241 dvss.n13 13.8526
R11510 dvss.n244 dvss.n9 13.8526
R11511 dvss.n221 dvss.n219 13.7605
R11512 dvss.n117 dvss.n116 13.6894
R11513 dvss.n75 dvss.n74 13.6894
R11514 dvss.n25 dvss.n24 13.5019
R11515 dvss.n223 dvss.n216 13.4405
R11516 dvss.n4141 dvss.n4140 13.4405
R11517 dvss.n4022 dvss.n4020 13.3
R11518 dvss.n4135 dvss.n4 13.2077
R11519 dvss.n3723 dvss.t10 13.1192
R11520 dvss.t359 dvss.n3649 13.1192
R11521 dvss.t321 dvss.n2203 13.1192
R11522 dvss.t52 dvss.n2178 13.1192
R11523 dvss.n2150 dvss.t443 13.1192
R11524 dvss.t317 dvss.n1991 13.1192
R11525 dvss.n1601 dvss.t648 13.1192
R11526 dvss.t349 dvss.n1516 13.1192
R11527 dvss.n1190 dvss.t155 13.1192
R11528 dvss.n211 dvss.n180 12.6405
R11529 dvss.n215 dvss.n182 12.6405
R11530 dvss.n3766 dvss.n3738 12.5222
R11531 dvss.n3687 dvss.n478 12.5222
R11532 dvss.n3009 dvss.n2126 12.5222
R11533 dvss.n3059 dvss.n2095 12.5222
R11534 dvss.n3109 dvss.n2064 12.5222
R11535 dvss.n2029 dvss.n714 12.5222
R11536 dvss.n1631 dvss.n1589 12.5222
R11537 dvss.n1554 dvss.n823 12.5222
R11538 dvss.n1158 dvss.n1157 12.5222
R11539 dvss.n3951 dvss.n3950 12.5222
R11540 dvss.n3886 dvss.n380 12.5222
R11541 dvss.n3485 dvss.n3482 12.5222
R11542 dvss.n3374 dvss.n3371 12.5222
R11543 dvss.n3253 dvss.n3250 12.5222
R11544 dvss.n1923 dvss.n1845 12.5222
R11545 dvss.n1775 dvss.n1772 12.5222
R11546 dvss.n1448 dvss.n1370 12.5222
R11547 dvss.n1300 dvss.n1297 12.5222
R11548 dvss.n194 dvss.n193 12.3205
R11549 dvss.n1006 dvss.n1005 12.2361
R11550 dvss.n2869 dvss.n2406 12.2361
R11551 dvss.n1087 dvss.n1085 12.1422
R11552 dvss.n1000 dvss.n999 12.1422
R11553 dvss.n3833 dvss.t141 11.3663
R11554 dvss.n3581 dvss.t475 11.3663
R11555 dvss.n3465 dvss.t192 11.3663
R11556 dvss.n3349 dvss.t22 11.3663
R11557 dvss.n3233 dvss.t632 11.3663
R11558 dvss.n1890 dvss.t464 11.3663
R11559 dvss.n1755 dvss.t673 11.3663
R11560 dvss.n1415 dvss.t505 11.3663
R11561 dvss.n1280 dvss.t418 11.3663
R11562 dvss.t0 dvss.t248 11.3596
R11563 dvss.n132 dvss.n131 11.2005
R11564 dvss.n87 dvss.n62 11.2005
R11565 dvss.n40 dvss.n39 11.0471
R11566 dvss.t248 dvss.t266 11.0256
R11567 dvss.n122 dvss.n121 10.8449
R11568 dvss.n79 dvss.n78 10.8449
R11569 dvss.n4136 dvss.n4135 10.7826
R11570 dvss.n30 dvss.n29 10.6964
R11571 dvss.n3713 dvss.t5 10.6405
R11572 dvss.n3713 dvss.t7 10.6405
R11573 dvss.n3706 dvss.t11 10.6405
R11574 dvss.n3706 dvss.t3 10.6405
R11575 dvss.n485 dvss.t364 10.6405
R11576 dvss.n485 dvss.t366 10.6405
R11577 dvss.n494 dvss.t360 10.6405
R11578 dvss.n494 dvss.t362 10.6405
R11579 dvss.n2117 dvss.t326 10.6405
R11580 dvss.n2117 dvss.t328 10.6405
R11581 dvss.n2111 dvss.t322 10.6405
R11582 dvss.n2111 dvss.t324 10.6405
R11583 dvss.n2086 dvss.t57 10.6405
R11584 dvss.n2086 dvss.t59 10.6405
R11585 dvss.n2080 dvss.t53 10.6405
R11586 dvss.n2080 dvss.t55 10.6405
R11587 dvss.n2055 dvss.t442 10.6405
R11588 dvss.n2055 dvss.t440 10.6405
R11589 dvss.n2048 dvss.t444 10.6405
R11590 dvss.n2048 dvss.t446 10.6405
R11591 dvss.n721 dvss.t314 10.6405
R11592 dvss.n721 dvss.t320 10.6405
R11593 dvss.n730 dvss.t318 10.6405
R11594 dvss.n730 dvss.t316 10.6405
R11595 dvss.n1580 dvss.t645 10.6405
R11596 dvss.n1580 dvss.t643 10.6405
R11597 dvss.n1573 dvss.t649 10.6405
R11598 dvss.n1573 dvss.t647 10.6405
R11599 dvss.n830 dvss.t348 10.6405
R11600 dvss.n830 dvss.t354 10.6405
R11601 dvss.n839 dvss.t350 10.6405
R11602 dvss.n839 dvss.t346 10.6405
R11603 dvss.n1136 dvss.t154 10.6405
R11604 dvss.n1136 dvss.t158 10.6405
R11605 dvss.n1128 dvss.t156 10.6405
R11606 dvss.n1128 dvss.t150 10.6405
R11607 dvss.n413 dvss.t140 10.6405
R11608 dvss.n413 dvss.t142 10.6405
R11609 dvss.n411 dvss.t136 10.6405
R11610 dvss.n411 dvss.t138 10.6405
R11611 dvss.n3534 dvss.t474 10.6405
R11612 dvss.n3534 dvss.t476 10.6405
R11613 dvss.n3532 dvss.t470 10.6405
R11614 dvss.n3532 dvss.t472 10.6405
R11615 dvss.n3452 dvss.t191 10.6405
R11616 dvss.n3452 dvss.t193 10.6405
R11617 dvss.n3432 dvss.t187 10.6405
R11618 dvss.n3432 dvss.t189 10.6405
R11619 dvss.n3334 dvss.t21 10.6405
R11620 dvss.n3334 dvss.t23 10.6405
R11621 dvss.n616 dvss.t17 10.6405
R11622 dvss.n616 dvss.t19 10.6405
R11623 dvss.n3220 dvss.t635 10.6405
R11624 dvss.n3220 dvss.t633 10.6405
R11625 dvss.n3206 dvss.t637 10.6405
R11626 dvss.n3206 dvss.t639 10.6405
R11627 dvss.n1824 dvss.t459 10.6405
R11628 dvss.n1824 dvss.t465 10.6405
R11629 dvss.n1822 dvss.t463 10.6405
R11630 dvss.n1822 dvss.t461 10.6405
R11631 dvss.n1742 dvss.t676 10.6405
R11632 dvss.n1742 dvss.t674 10.6405
R11633 dvss.n1728 dvss.t680 10.6405
R11634 dvss.n1728 dvss.t678 10.6405
R11635 dvss.n1349 dvss.t510 10.6405
R11636 dvss.n1349 dvss.t506 10.6405
R11637 dvss.n1347 dvss.t512 10.6405
R11638 dvss.n1347 dvss.t508 10.6405
R11639 dvss.n1267 dvss.t425 10.6405
R11640 dvss.n1267 dvss.t419 10.6405
R11641 dvss.n1253 dvss.t427 10.6405
R11642 dvss.n1253 dvss.t421 10.6405
R11643 dvss.n334 dvss.t209 10.6405
R11644 dvss.n334 dvss.t213 10.6405
R11645 dvss.n337 dvss.t207 10.6405
R11646 dvss.n337 dvss.t215 10.6405
R11647 dvss.n385 dvss.t128 10.6405
R11648 dvss.n385 dvss.t124 10.6405
R11649 dvss.n3880 dvss.t132 10.6405
R11650 dvss.n3880 dvss.t134 10.6405
R11651 dvss.n519 dvss.t33 10.6405
R11652 dvss.n519 dvss.t27 10.6405
R11653 dvss.n522 dvss.t35 10.6405
R11654 dvss.n522 dvss.t29 10.6405
R11655 dvss.n582 dvss.t39 10.6405
R11656 dvss.n582 dvss.t41 10.6405
R11657 dvss.n585 dvss.t47 10.6405
R11658 dvss.n585 dvss.t43 10.6405
R11659 dvss.n645 dvss.t302 10.6405
R11660 dvss.n645 dvss.t300 10.6405
R11661 dvss.n648 dvss.t298 10.6405
R11662 dvss.n648 dvss.t296 10.6405
R11663 dvss.n1840 dvss.t574 10.6405
R11664 dvss.n1840 dvss.t566 10.6405
R11665 dvss.n1917 dvss.t572 10.6405
R11666 dvss.n1917 dvss.t570 10.6405
R11667 dvss.n754 dvss.t290 10.6405
R11668 dvss.n754 dvss.t288 10.6405
R11669 dvss.n757 dvss.t286 10.6405
R11670 dvss.n757 dvss.t280 10.6405
R11671 dvss.n1365 dvss.t593 10.6405
R11672 dvss.n1365 dvss.t591 10.6405
R11673 dvss.n1442 dvss.t589 10.6405
R11674 dvss.n1442 dvss.t587 10.6405
R11675 dvss.n863 dvss.t344 10.6405
R11676 dvss.n863 dvss.t342 10.6405
R11677 dvss.n866 dvss.t340 10.6405
R11678 dvss.n866 dvss.t338 10.6405
R11679 dvss.n4082 dvss.t662 10.6405
R11680 dvss.n4082 dvss.t666 10.6405
R11681 dvss.n4074 dvss.t660 10.6405
R11682 dvss.n4074 dvss.t668 10.6405
R11683 dvss.n4115 dvss.t179 10.6405
R11684 dvss.n4115 dvss.t175 10.6405
R11685 dvss.n269 dvss.t183 10.6405
R11686 dvss.n269 dvss.t185 10.6405
R11687 dvss.n2288 dvss.t261 10.6405
R11688 dvss.n2288 dvss.t255 10.6405
R11689 dvss.n2214 dvss.t263 10.6405
R11690 dvss.n2214 dvss.t257 10.6405
R11691 dvss.n2308 dvss.t110 10.6405
R11692 dvss.n2308 dvss.t112 10.6405
R11693 dvss.n2311 dvss.t118 10.6405
R11694 dvss.n2311 dvss.t114 10.6405
R11695 dvss.n2644 dvss.t544 10.6405
R11696 dvss.n2644 dvss.t543 10.6405
R11697 dvss.n2636 dvss.t542 10.6405
R11698 dvss.n2636 dvss.t541 10.6405
R11699 dvss.n2691 dvss.t581 10.6405
R11700 dvss.n2691 dvss.t577 10.6405
R11701 dvss.n2683 dvss.t580 10.6405
R11702 dvss.n2683 dvss.t579 10.6405
R11703 dvss.n2738 dvss.t533 10.6405
R11704 dvss.n2738 dvss.t532 10.6405
R11705 dvss.n2730 dvss.t531 10.6405
R11706 dvss.n2730 dvss.t527 10.6405
R11707 dvss.n2785 dvss.t205 10.6405
R11708 dvss.n2785 dvss.t204 10.6405
R11709 dvss.n2777 dvss.t203 10.6405
R11710 dvss.n2777 dvss.t202 10.6405
R11711 dvss.n2832 dvss.t245 10.6405
R11712 dvss.n2832 dvss.t244 10.6405
R11713 dvss.n2824 dvss.t243 10.6405
R11714 dvss.n2824 dvss.t242 10.6405
R11715 dvss.n3793 dvss.n3792 10.64
R11716 dvss.n3643 dvss.n495 10.64
R11717 dvss.n3036 dvss.n3035 10.64
R11718 dvss.n3086 dvss.n3085 10.64
R11719 dvss.n3136 dvss.n3135 10.64
R11720 dvss.n1985 dvss.n731 10.64
R11721 dvss.n1658 dvss.n1657 10.64
R11722 dvss.n1510 dvss.n840 10.64
R11723 dvss.n1129 dvss.n1127 10.64
R11724 dvss.n412 dvss.n410 10.64
R11725 dvss.n3533 dvss.n3531 10.64
R11726 dvss.n3437 dvss.n3436 10.64
R11727 dvss.n625 dvss.n617 10.64
R11728 dvss.n3207 dvss.n3205 10.64
R11729 dvss.n1823 dvss.n1821 10.64
R11730 dvss.n1729 dvss.n1727 10.64
R11731 dvss.n1348 dvss.n1346 10.64
R11732 dvss.n1254 dvss.n1252 10.64
R11733 dvss.n4027 dvss.n4009 10.6369
R11734 dvss.n4031 dvss.n4009 10.6369
R11735 dvss.n4030 dvss.n4029 10.6369
R11736 dvss.n4031 dvss.n4030 10.6369
R11737 dvss.n4007 dvss.n4006 10.6369
R11738 dvss.n4010 dvss.n4007 10.6369
R11739 dvss.n4036 dvss.n3993 10.6369
R11740 dvss.n4010 dvss.n3993 10.6369
R11741 dvss.n153 dvss.n152 10.3672
R11742 dvss.n155 dvss.n97 10.3672
R11743 dvss.n256 dvss.n255 10.3526
R11744 dvss.n209 dvss.n208 10.0805
R11745 dvss.t606 dvss.n234 10.0615
R11746 dvss.n199 dvss.n198 9.7605
R11747 dvss.n2887 dvss 9.31486
R11748 dvss.n1229 dvss 9.30735
R11749 dvss.n963 dvss.n914 9.30085
R11750 dvss.n1007 dvss.n1006 9.3005
R11751 dvss.n1006 dvss.n1002 9.3005
R11752 dvss.n1024 dvss.n1019 9.3005
R11753 dvss.n1025 dvss.n1024 9.3005
R11754 dvss.n1243 dvss.n1242 9.3005
R11755 dvss.n1242 dvss.n1239 9.3005
R11756 dvss.n1324 dvss.n860 9.3005
R11757 dvss.n1325 dvss.n1324 9.3005
R11758 dvss.n1322 dvss.n865 9.3005
R11759 dvss.n1322 dvss.n1321 9.3005
R11760 dvss.n1292 dvss.n864 9.3005
R11761 dvss.n881 dvss.n864 9.3005
R11762 dvss.n1476 dvss.n1475 9.3005
R11763 dvss.n1477 dvss.n1476 9.3005
R11764 dvss.n1682 dvss.n1681 9.3005
R11765 dvss.n1681 dvss.n1680 9.3005
R11766 dvss.n1445 dvss.n1444 9.3005
R11767 dvss.n1444 dvss.n1443 9.3005
R11768 dvss.n1367 dvss.n1366 9.3005
R11769 dvss.n1366 dvss.n1359 9.3005
R11770 dvss.n1718 dvss.n1717 9.3005
R11771 dvss.n1717 dvss.n1714 9.3005
R11772 dvss.n1799 dvss.n751 9.3005
R11773 dvss.n1800 dvss.n1799 9.3005
R11774 dvss.n1797 dvss.n756 9.3005
R11775 dvss.n1797 dvss.n1796 9.3005
R11776 dvss.n1767 dvss.n755 9.3005
R11777 dvss.n772 dvss.n755 9.3005
R11778 dvss.n1951 dvss.n1950 9.3005
R11779 dvss.n1952 dvss.n1951 9.3005
R11780 dvss.n3160 dvss.n3159 9.3005
R11781 dvss.n3159 dvss.n3158 9.3005
R11782 dvss.n1920 dvss.n1919 9.3005
R11783 dvss.n1919 dvss.n1918 9.3005
R11784 dvss.n1842 dvss.n1841 9.3005
R11785 dvss.n1841 dvss.n1834 9.3005
R11786 dvss.n3196 dvss.n3195 9.3005
R11787 dvss.n3195 dvss.n3192 9.3005
R11788 dvss.n3278 dvss.n641 9.3005
R11789 dvss.n3279 dvss.n3278 9.3005
R11790 dvss.n3276 dvss.n647 9.3005
R11791 dvss.n3276 dvss.n3275 9.3005
R11792 dvss.n3245 dvss.n646 9.3005
R11793 dvss.n663 dvss.n646 9.3005
R11794 dvss.n3315 dvss.n3314 9.3005
R11795 dvss.n3314 dvss.n3311 9.3005
R11796 dvss.n3395 dvss.n579 9.3005
R11797 dvss.n3396 dvss.n3395 9.3005
R11798 dvss.n3393 dvss.n584 9.3005
R11799 dvss.n3393 dvss.n3392 9.3005
R11800 dvss.n3361 dvss.n583 9.3005
R11801 dvss.n603 dvss.n583 9.3005
R11802 dvss.n3428 dvss.n3427 9.3005
R11803 dvss.n3427 dvss.n3424 9.3005
R11804 dvss.n3509 dvss.n516 9.3005
R11805 dvss.n3510 dvss.n3509 9.3005
R11806 dvss.n3507 dvss.n521 9.3005
R11807 dvss.n3507 dvss.n3506 9.3005
R11808 dvss.n3477 dvss.n520 9.3005
R11809 dvss.n537 dvss.n520 9.3005
R11810 dvss.n3609 dvss.n3608 9.3005
R11811 dvss.n3610 dvss.n3609 9.3005
R11812 dvss.n3878 dvss.n3877 9.3005
R11813 dvss.n3878 dvss.n387 9.3005
R11814 dvss.n3883 dvss.n3882 9.3005
R11815 dvss.n3882 dvss.n3881 9.3005
R11816 dvss.n386 dvss.n384 9.3005
R11817 dvss.n3587 dvss.n386 9.3005
R11818 dvss.n3865 dvss.n3864 9.3005
R11819 dvss.n3866 dvss.n3865 9.3005
R11820 dvss.n3960 dvss.n322 9.3005
R11821 dvss.n3961 dvss.n3960 9.3005
R11822 dvss.n3958 dvss.n336 9.3005
R11823 dvss.n3958 dvss.n3957 9.3005
R11824 dvss.n3936 dvss.n335 9.3005
R11825 dvss.n3843 dvss.n335 9.3005
R11826 dvss.n986 dvss.n985 9.3005
R11827 dvss.n985 dvss.n984 9.3005
R11828 dvss.n1028 dvss.n1027 9.3005
R11829 dvss.n1027 dvss.n1026 9.3005
R11830 dvss.n1299 dvss.n868 9.3005
R11831 dvss.n1297 dvss.n1296 9.3005
R11832 dvss.n1290 dvss.n1289 9.3005
R11833 dvss.n1256 dvss.n1255 9.3005
R11834 dvss.n1266 dvss.n1265 9.3005
R11835 dvss.n1271 dvss.n1270 9.3005
R11836 dvss.n1291 dvss.n1290 9.3005
R11837 dvss.n1447 dvss.n1446 9.3005
R11838 dvss.n1441 dvss.n1370 9.3005
R11839 dvss.n1460 dvss.n1459 9.3005
R11840 dvss.n1470 dvss.n1469 9.3005
R11841 dvss.n1467 dvss.n1466 9.3005
R11842 dvss.n1457 dvss.n1456 9.3005
R11843 dvss.n1459 dvss.n1455 9.3005
R11844 dvss.n1774 dvss.n759 9.3005
R11845 dvss.n1772 dvss.n1771 9.3005
R11846 dvss.n1765 dvss.n1764 9.3005
R11847 dvss.n1731 dvss.n1730 9.3005
R11848 dvss.n1741 dvss.n1740 9.3005
R11849 dvss.n1746 dvss.n1745 9.3005
R11850 dvss.n1766 dvss.n1765 9.3005
R11851 dvss.n1922 dvss.n1921 9.3005
R11852 dvss.n1916 dvss.n1845 9.3005
R11853 dvss.n1935 dvss.n1934 9.3005
R11854 dvss.n1945 dvss.n1944 9.3005
R11855 dvss.n1942 dvss.n1941 9.3005
R11856 dvss.n1932 dvss.n1931 9.3005
R11857 dvss.n1934 dvss.n1930 9.3005
R11858 dvss.n3252 dvss.n650 9.3005
R11859 dvss.n3250 dvss.n3249 9.3005
R11860 dvss.n3243 dvss.n3242 9.3005
R11861 dvss.n3209 dvss.n3208 9.3005
R11862 dvss.n3219 dvss.n3218 9.3005
R11863 dvss.n3224 dvss.n3223 9.3005
R11864 dvss.n3244 dvss.n3243 9.3005
R11865 dvss.n3373 dvss.n587 9.3005
R11866 dvss.n3371 dvss.n3370 9.3005
R11867 dvss.n3359 dvss.n3358 9.3005
R11868 dvss.n3332 dvss.n3331 9.3005
R11869 dvss.n3341 dvss.n3340 9.3005
R11870 dvss.n3338 dvss.n3337 9.3005
R11871 dvss.n3360 dvss.n3359 9.3005
R11872 dvss.n3484 dvss.n524 9.3005
R11873 dvss.n3482 dvss.n3481 9.3005
R11874 dvss.n3475 dvss.n3474 9.3005
R11875 dvss.n3435 dvss.n3434 9.3005
R11876 dvss.n3451 dvss.n3450 9.3005
R11877 dvss.n3456 dvss.n3455 9.3005
R11878 dvss.n3476 dvss.n3475 9.3005
R11879 dvss.n3885 dvss.n3884 9.3005
R11880 dvss.n383 dvss.n380 9.3005
R11881 dvss.n3593 dvss.n3592 9.3005
R11882 dvss.n3603 dvss.n3602 9.3005
R11883 dvss.n3600 dvss.n3599 9.3005
R11884 dvss.n3590 dvss.n3589 9.3005
R11885 dvss.n3592 dvss.n3588 9.3005
R11886 dvss.n3949 dvss.n339 9.3005
R11887 dvss.n3952 dvss.n3951 9.3005
R11888 dvss.n3849 dvss.n3848 9.3005
R11889 dvss.n3859 dvss.n3858 9.3005
R11890 dvss.n3856 dvss.n3855 9.3005
R11891 dvss.n3846 dvss.n3845 9.3005
R11892 dvss.n3848 dvss.n3844 9.3005
R11893 dvss.n1000 dvss.n997 9.3005
R11894 dvss.n1001 dvss.n1000 9.3005
R11895 dvss.n1076 dvss.n1075 9.3005
R11896 dvss.n1075 dvss.n1074 9.3005
R11897 dvss.n1101 dvss.n1100 9.3005
R11898 dvss.n1100 dvss.n1099 9.3005
R11899 dvss.n1156 dvss.n1155 9.3005
R11900 dvss.n1159 dvss.n1158 9.3005
R11901 dvss.n1143 dvss.n1142 9.3005
R11902 dvss.n1131 dvss.n1130 9.3005
R11903 dvss.n1135 dvss.n1134 9.3005
R11904 dvss.n1139 dvss.n1138 9.3005
R11905 dvss.n1144 dvss.n1143 9.3005
R11906 dvss.n1556 dvss.n1555 9.3005
R11907 dvss.n823 dvss.n822 9.3005
R11908 dvss.n1540 dvss.n828 9.3005
R11909 dvss.n1523 dvss.n1522 9.3005
R11910 dvss.n1526 dvss.n1525 9.3005
R11911 dvss.n1538 dvss.n1537 9.3005
R11912 dvss.n1541 dvss.n1540 9.3005
R11913 dvss.n1630 dvss.n1629 9.3005
R11914 dvss.n1628 dvss.n1589 9.3005
R11915 dvss.n1641 dvss.n1640 9.3005
R11916 dvss.n1656 dvss.n1655 9.3005
R11917 dvss.n1650 dvss.n1649 9.3005
R11918 dvss.n1647 dvss.n1646 9.3005
R11919 dvss.n1640 dvss.n1638 9.3005
R11920 dvss.n2031 dvss.n2030 9.3005
R11921 dvss.n714 dvss.n713 9.3005
R11922 dvss.n2015 dvss.n719 9.3005
R11923 dvss.n1998 dvss.n1997 9.3005
R11924 dvss.n2001 dvss.n2000 9.3005
R11925 dvss.n2013 dvss.n2012 9.3005
R11926 dvss.n2016 dvss.n2015 9.3005
R11927 dvss.n3108 dvss.n3107 9.3005
R11928 dvss.n3106 dvss.n2064 9.3005
R11929 dvss.n3119 dvss.n3118 9.3005
R11930 dvss.n3134 dvss.n3133 9.3005
R11931 dvss.n3128 dvss.n3127 9.3005
R11932 dvss.n3125 dvss.n3124 9.3005
R11933 dvss.n3118 dvss.n3116 9.3005
R11934 dvss.n3058 dvss.n3057 9.3005
R11935 dvss.n3056 dvss.n2095 9.3005
R11936 dvss.n3069 dvss.n3068 9.3005
R11937 dvss.n3084 dvss.n3083 9.3005
R11938 dvss.n3078 dvss.n3077 9.3005
R11939 dvss.n3075 dvss.n3074 9.3005
R11940 dvss.n3068 dvss.n3066 9.3005
R11941 dvss.n3008 dvss.n3007 9.3005
R11942 dvss.n3006 dvss.n2126 9.3005
R11943 dvss.n3019 dvss.n3018 9.3005
R11944 dvss.n3034 dvss.n3033 9.3005
R11945 dvss.n3028 dvss.n3027 9.3005
R11946 dvss.n3025 dvss.n3024 9.3005
R11947 dvss.n3018 dvss.n3016 9.3005
R11948 dvss.n3689 dvss.n3688 9.3005
R11949 dvss.n478 dvss.n477 9.3005
R11950 dvss.n3673 dvss.n483 9.3005
R11951 dvss.n3656 dvss.n3655 9.3005
R11952 dvss.n3659 dvss.n3658 9.3005
R11953 dvss.n3671 dvss.n3670 9.3005
R11954 dvss.n3674 dvss.n3673 9.3005
R11955 dvss.n3765 dvss.n3764 9.3005
R11956 dvss.n3763 dvss.n3738 9.3005
R11957 dvss.n3776 dvss.n3775 9.3005
R11958 dvss.n3791 dvss.n3790 9.3005
R11959 dvss.n3785 dvss.n3784 9.3005
R11960 dvss.n3782 dvss.n3781 9.3005
R11961 dvss.n3775 dvss.n3773 9.3005
R11962 dvss.n1088 dvss.n1087 9.3005
R11963 dvss.n1087 dvss.n1086 9.3005
R11964 dvss.n1228 dvss.n1059 9.3005
R11965 dvss.n1227 dvss.n1060 9.3005
R11966 dvss.n1065 dvss.n1061 9.3005
R11967 dvss.n1221 dvss.n1066 9.3005
R11968 dvss.n1220 dvss.n1067 9.3005
R11969 dvss.n1219 dvss.n1068 9.3005
R11970 dvss.n1073 dvss.n1069 9.3005
R11971 dvss.n1212 dvss.n1077 9.3005
R11972 dvss.n1211 dvss.n1078 9.3005
R11973 dvss.n1210 dvss.n1079 9.3005
R11974 dvss.n1089 dvss.n1080 9.3005
R11975 dvss.n1204 dvss.n1090 9.3005
R11976 dvss.n1203 dvss.n1091 9.3005
R11977 dvss.n1202 dvss.n1092 9.3005
R11978 dvss.n1102 dvss.n1093 9.3005
R11979 dvss.n1196 dvss.n1103 9.3005
R11980 dvss.n1195 dvss.n1104 9.3005
R11981 dvss.n1194 dvss.n1105 9.3005
R11982 dvss.n1109 dvss.n1106 9.3005
R11983 dvss.n1188 dvss.n1110 9.3005
R11984 dvss.n1187 dvss.n1111 9.3005
R11985 dvss.n1186 dvss.n1112 9.3005
R11986 dvss.n1133 dvss.n1113 9.3005
R11987 dvss.n1180 dvss.n1117 9.3005
R11988 dvss.n1179 dvss.n1118 9.3005
R11989 dvss.n1178 dvss.n1119 9.3005
R11990 dvss.n1141 dvss.n1120 9.3005
R11991 dvss.n1172 dvss.n1145 9.3005
R11992 dvss.n1171 dvss.n1146 9.3005
R11993 dvss.n1170 dvss.n1147 9.3005
R11994 dvss.n1154 dvss.n1148 9.3005
R11995 dvss.n1164 dvss.n1160 9.3005
R11996 dvss.n1163 dvss.n1162 9.3005
R11997 dvss.n1161 dvss.n850 9.3005
R11998 dvss.n1497 dvss.n1496 9.3005
R11999 dvss.n1498 dvss.n849 9.3005
R12000 dvss.n1501 dvss.n1500 9.3005
R12001 dvss.n1499 dvss.n846 9.3005
R12002 dvss.n1508 dvss.n1507 9.3005
R12003 dvss.n1509 dvss.n845 9.3005
R12004 dvss.n1513 dvss.n1512 9.3005
R12005 dvss.n1511 dvss.n841 9.3005
R12006 dvss.n1520 dvss.n1519 9.3005
R12007 dvss.n1521 dvss.n837 9.3005
R12008 dvss.n1528 dvss.n1527 9.3005
R12009 dvss.n838 dvss.n833 9.3005
R12010 dvss.n1536 dvss.n1535 9.3005
R12011 dvss.n832 dvss.n827 9.3005
R12012 dvss.n1543 dvss.n1542 9.3005
R12013 dvss.n829 dvss.n824 9.3005
R12014 dvss.n1551 dvss.n1550 9.3005
R12015 dvss.n1552 dvss.n819 9.3005
R12016 dvss.n1558 dvss.n1557 9.3005
R12017 dvss.n821 dvss.n816 9.3005
R12018 dvss.n1565 dvss.n1564 9.3005
R12019 dvss.n1566 dvss.n814 9.3005
R12020 dvss.n1671 dvss.n1670 9.3005
R12021 dvss.n1669 dvss.n815 9.3005
R12022 dvss.n1668 dvss.n1667 9.3005
R12023 dvss.n1666 dvss.n1665 9.3005
R12024 dvss.n1664 dvss.n1569 9.3005
R12025 dvss.n1663 dvss.n1662 9.3005
R12026 dvss.n1661 dvss.n1660 9.3005
R12027 dvss.n1659 dvss.n1572 9.3005
R12028 dvss.n1575 dvss.n1574 9.3005
R12029 dvss.n1654 dvss.n1653 9.3005
R12030 dvss.n1652 dvss.n1651 9.3005
R12031 dvss.n1581 dvss.n1578 9.3005
R12032 dvss.n1645 dvss.n1644 9.3005
R12033 dvss.n1643 dvss.n1642 9.3005
R12034 dvss.n1585 dvss.n1584 9.3005
R12035 dvss.n1637 dvss.n1636 9.3005
R12036 dvss.n1635 dvss.n1634 9.3005
R12037 dvss.n1633 dvss.n1588 9.3005
R12038 dvss.n1592 dvss.n1591 9.3005
R12039 dvss.n1627 dvss.n1626 9.3005
R12040 dvss.n1625 dvss.n1624 9.3005
R12041 dvss.n1623 dvss.n741 9.3005
R12042 dvss.n1972 dvss.n1971 9.3005
R12043 dvss.n1973 dvss.n740 9.3005
R12044 dvss.n1976 dvss.n1975 9.3005
R12045 dvss.n1974 dvss.n737 9.3005
R12046 dvss.n1983 dvss.n1982 9.3005
R12047 dvss.n1984 dvss.n736 9.3005
R12048 dvss.n1988 dvss.n1987 9.3005
R12049 dvss.n1986 dvss.n732 9.3005
R12050 dvss.n1995 dvss.n1994 9.3005
R12051 dvss.n1996 dvss.n728 9.3005
R12052 dvss.n2003 dvss.n2002 9.3005
R12053 dvss.n729 dvss.n724 9.3005
R12054 dvss.n2011 dvss.n2010 9.3005
R12055 dvss.n723 dvss.n718 9.3005
R12056 dvss.n2018 dvss.n2017 9.3005
R12057 dvss.n720 dvss.n715 9.3005
R12058 dvss.n2026 dvss.n2025 9.3005
R12059 dvss.n2027 dvss.n710 9.3005
R12060 dvss.n2033 dvss.n2032 9.3005
R12061 dvss.n712 dvss.n707 9.3005
R12062 dvss.n2040 dvss.n2039 9.3005
R12063 dvss.n2041 dvss.n705 9.3005
R12064 dvss.n3149 dvss.n3148 9.3005
R12065 dvss.n3147 dvss.n706 9.3005
R12066 dvss.n3146 dvss.n3145 9.3005
R12067 dvss.n3144 dvss.n3143 9.3005
R12068 dvss.n3142 dvss.n2044 9.3005
R12069 dvss.n3141 dvss.n3140 9.3005
R12070 dvss.n3139 dvss.n3138 9.3005
R12071 dvss.n3137 dvss.n2047 9.3005
R12072 dvss.n2050 dvss.n2049 9.3005
R12073 dvss.n3132 dvss.n3131 9.3005
R12074 dvss.n3130 dvss.n3129 9.3005
R12075 dvss.n2056 dvss.n2053 9.3005
R12076 dvss.n3123 dvss.n3122 9.3005
R12077 dvss.n3121 dvss.n3120 9.3005
R12078 dvss.n2060 dvss.n2059 9.3005
R12079 dvss.n3115 dvss.n3114 9.3005
R12080 dvss.n3113 dvss.n3112 9.3005
R12081 dvss.n3111 dvss.n2063 9.3005
R12082 dvss.n2067 dvss.n2066 9.3005
R12083 dvss.n3105 dvss.n3104 9.3005
R12084 dvss.n3103 dvss.n3102 9.3005
R12085 dvss.n3101 dvss.n2070 9.3005
R12086 dvss.n3100 dvss.n3099 9.3005
R12087 dvss.n3098 dvss.n3097 9.3005
R12088 dvss.n3096 dvss.n2073 9.3005
R12089 dvss.n3095 dvss.n3094 9.3005
R12090 dvss.n3093 dvss.n3092 9.3005
R12091 dvss.n3091 dvss.n2076 9.3005
R12092 dvss.n3090 dvss.n3089 9.3005
R12093 dvss.n3088 dvss.n3087 9.3005
R12094 dvss.n2081 dvss.n2079 9.3005
R12095 dvss.n3082 dvss.n3081 9.3005
R12096 dvss.n3080 dvss.n3079 9.3005
R12097 dvss.n2087 dvss.n2084 9.3005
R12098 dvss.n3073 dvss.n3072 9.3005
R12099 dvss.n3071 dvss.n3070 9.3005
R12100 dvss.n2091 dvss.n2090 9.3005
R12101 dvss.n3065 dvss.n3064 9.3005
R12102 dvss.n3063 dvss.n3062 9.3005
R12103 dvss.n3061 dvss.n2094 9.3005
R12104 dvss.n2098 dvss.n2097 9.3005
R12105 dvss.n3055 dvss.n3054 9.3005
R12106 dvss.n3053 dvss.n3052 9.3005
R12107 dvss.n3051 dvss.n2101 9.3005
R12108 dvss.n3050 dvss.n3049 9.3005
R12109 dvss.n3048 dvss.n3047 9.3005
R12110 dvss.n3046 dvss.n2104 9.3005
R12111 dvss.n3045 dvss.n3044 9.3005
R12112 dvss.n3043 dvss.n3042 9.3005
R12113 dvss.n3041 dvss.n2107 9.3005
R12114 dvss.n3040 dvss.n3039 9.3005
R12115 dvss.n3038 dvss.n3037 9.3005
R12116 dvss.n2112 dvss.n2110 9.3005
R12117 dvss.n3032 dvss.n3031 9.3005
R12118 dvss.n3030 dvss.n3029 9.3005
R12119 dvss.n2118 dvss.n2115 9.3005
R12120 dvss.n3023 dvss.n3022 9.3005
R12121 dvss.n3021 dvss.n3020 9.3005
R12122 dvss.n2122 dvss.n2121 9.3005
R12123 dvss.n3015 dvss.n3014 9.3005
R12124 dvss.n3013 dvss.n3012 9.3005
R12125 dvss.n3011 dvss.n2125 9.3005
R12126 dvss.n2129 dvss.n2128 9.3005
R12127 dvss.n3005 dvss.n3004 9.3005
R12128 dvss.n3003 dvss.n3002 9.3005
R12129 dvss.n3001 dvss.n505 9.3005
R12130 dvss.n3630 dvss.n3629 9.3005
R12131 dvss.n3631 dvss.n504 9.3005
R12132 dvss.n3634 dvss.n3633 9.3005
R12133 dvss.n3632 dvss.n501 9.3005
R12134 dvss.n3641 dvss.n3640 9.3005
R12135 dvss.n3642 dvss.n500 9.3005
R12136 dvss.n3646 dvss.n3645 9.3005
R12137 dvss.n3644 dvss.n496 9.3005
R12138 dvss.n3653 dvss.n3652 9.3005
R12139 dvss.n3654 dvss.n492 9.3005
R12140 dvss.n3661 dvss.n3660 9.3005
R12141 dvss.n493 dvss.n488 9.3005
R12142 dvss.n3669 dvss.n3668 9.3005
R12143 dvss.n487 dvss.n482 9.3005
R12144 dvss.n3676 dvss.n3675 9.3005
R12145 dvss.n484 dvss.n479 9.3005
R12146 dvss.n3684 dvss.n3683 9.3005
R12147 dvss.n3685 dvss.n474 9.3005
R12148 dvss.n3691 dvss.n3690 9.3005
R12149 dvss.n476 dvss.n471 9.3005
R12150 dvss.n3698 dvss.n3697 9.3005
R12151 dvss.n3699 dvss.n469 9.3005
R12152 dvss.n3806 dvss.n3805 9.3005
R12153 dvss.n3804 dvss.n470 9.3005
R12154 dvss.n3803 dvss.n3802 9.3005
R12155 dvss.n3801 dvss.n3800 9.3005
R12156 dvss.n3799 dvss.n3702 9.3005
R12157 dvss.n3798 dvss.n3797 9.3005
R12158 dvss.n3796 dvss.n3795 9.3005
R12159 dvss.n3794 dvss.n3705 9.3005
R12160 dvss.n3708 dvss.n3707 9.3005
R12161 dvss.n3789 dvss.n3788 9.3005
R12162 dvss.n3787 dvss.n3786 9.3005
R12163 dvss.n3714 dvss.n3711 9.3005
R12164 dvss.n3780 dvss.n3779 9.3005
R12165 dvss.n3778 dvss.n3777 9.3005
R12166 dvss.n3734 dvss.n3733 9.3005
R12167 dvss.n3772 dvss.n3771 9.3005
R12168 dvss.n3770 dvss.n3769 9.3005
R12169 dvss.n3768 dvss.n3737 9.3005
R12170 dvss.n3741 dvss.n3740 9.3005
R12171 dvss.n3762 dvss.n3761 9.3005
R12172 dvss.n3760 dvss.n3759 9.3005
R12173 dvss.n3758 dvss.n3756 9.3005
R12174 dvss.n3757 dvss.n311 9.3005
R12175 dvss.n4051 dvss.n4050 9.3005
R12176 dvss.n4049 dvss.n312 9.3005
R12177 dvss.n4048 dvss.n4047 9.3005
R12178 dvss.n962 dvss.n961 9.3005
R12179 dvss.n960 dvss.n959 9.3005
R12180 dvss.n970 dvss.n969 9.3005
R12181 dvss.n973 dvss.n972 9.3005
R12182 dvss.n975 dvss.n974 9.3005
R12183 dvss.n957 dvss.n956 9.3005
R12184 dvss.n983 dvss.n981 9.3005
R12185 dvss.n988 dvss.n987 9.3005
R12186 dvss.n990 dvss.n989 9.3005
R12187 dvss.n954 dvss.n953 9.3005
R12188 dvss.n1007 dvss.n996 9.3005
R12189 dvss.n1010 dvss.n1009 9.3005
R12190 dvss.n1012 dvss.n1011 9.3005
R12191 dvss.n935 dvss.n933 9.3005
R12192 dvss.n1018 dvss.n1017 9.3005
R12193 dvss.n939 dvss.n936 9.3005
R12194 dvss.n949 dvss.n948 9.3005
R12195 dvss.n1238 dvss.n902 9.3005
R12196 dvss.n901 dvss.n900 9.3005
R12197 dvss.n1245 dvss.n1244 9.3005
R12198 dvss.n1251 dvss.n896 9.3005
R12199 dvss.n1258 dvss.n1257 9.3005
R12200 dvss.n1264 dvss.n888 9.3005
R12201 dvss.n1273 dvss.n1272 9.3005
R12202 dvss.n1276 dvss.n1274 9.3005
R12203 dvss.n1275 dvss.n885 9.3005
R12204 dvss.n1288 dvss.n879 9.3005
R12205 dvss.n1294 dvss.n1293 9.3005
R12206 dvss.n1303 dvss.n1295 9.3005
R12207 dvss.n1302 dvss.n875 9.3005
R12208 dvss.n1320 dvss.n867 9.3005
R12209 dvss.n1317 dvss.n872 9.3005
R12210 dvss.n1316 dvss.n1315 9.3005
R12211 dvss.n1326 dvss.n858 9.3005
R12212 dvss.n1488 dvss.n1487 9.3005
R12213 dvss.n1484 dvss.n859 9.3005
R12214 dvss.n1483 dvss.n1330 9.3005
R12215 dvss.n1482 dvss.n1331 9.3005
R12216 dvss.n1479 dvss.n1335 9.3005
R12217 dvss.n1478 dvss.n1336 9.3005
R12218 dvss.n1401 dvss.n1339 9.3005
R12219 dvss.n1474 dvss.n1340 9.3005
R12220 dvss.n1471 dvss.n1345 9.3005
R12221 dvss.n1409 dvss.n1408 9.3005
R12222 dvss.n1411 dvss.n1410 9.3005
R12223 dvss.n1465 dvss.n1351 9.3005
R12224 dvss.n1462 dvss.n1356 9.3005
R12225 dvss.n1461 dvss.n1357 9.3005
R12226 dvss.n1378 dvss.n1358 9.3005
R12227 dvss.n1454 dvss.n1360 9.3005
R12228 dvss.n1451 dvss.n1368 9.3005
R12229 dvss.n1450 dvss.n1369 9.3005
R12230 dvss.n1377 dvss.n1372 9.3005
R12231 dvss.n1440 dvss.n1373 9.3005
R12232 dvss.n1437 dvss.n807 9.3005
R12233 dvss.n1679 dvss.n1678 9.3005
R12234 dvss.n1683 dvss.n802 9.3005
R12235 dvss.n1705 dvss.n1704 9.3005
R12236 dvss.n1701 dvss.n803 9.3005
R12237 dvss.n1700 dvss.n1692 9.3005
R12238 dvss.n1699 dvss.n1698 9.3005
R12239 dvss.n1713 dvss.n793 9.3005
R12240 dvss.n792 dvss.n791 9.3005
R12241 dvss.n1720 dvss.n1719 9.3005
R12242 dvss.n1726 dvss.n787 9.3005
R12243 dvss.n1733 dvss.n1732 9.3005
R12244 dvss.n1739 dvss.n779 9.3005
R12245 dvss.n1748 dvss.n1747 9.3005
R12246 dvss.n1751 dvss.n1749 9.3005
R12247 dvss.n1750 dvss.n776 9.3005
R12248 dvss.n1763 dvss.n770 9.3005
R12249 dvss.n1769 dvss.n1768 9.3005
R12250 dvss.n1778 dvss.n1770 9.3005
R12251 dvss.n1777 dvss.n766 9.3005
R12252 dvss.n1795 dvss.n758 9.3005
R12253 dvss.n1792 dvss.n763 9.3005
R12254 dvss.n1791 dvss.n1790 9.3005
R12255 dvss.n1801 dvss.n749 9.3005
R12256 dvss.n1963 dvss.n1962 9.3005
R12257 dvss.n1959 dvss.n750 9.3005
R12258 dvss.n1958 dvss.n1805 9.3005
R12259 dvss.n1957 dvss.n1806 9.3005
R12260 dvss.n1954 dvss.n1810 9.3005
R12261 dvss.n1953 dvss.n1811 9.3005
R12262 dvss.n1876 dvss.n1814 9.3005
R12263 dvss.n1949 dvss.n1815 9.3005
R12264 dvss.n1946 dvss.n1820 9.3005
R12265 dvss.n1884 dvss.n1883 9.3005
R12266 dvss.n1886 dvss.n1885 9.3005
R12267 dvss.n1940 dvss.n1826 9.3005
R12268 dvss.n1937 dvss.n1831 9.3005
R12269 dvss.n1936 dvss.n1832 9.3005
R12270 dvss.n1853 dvss.n1833 9.3005
R12271 dvss.n1929 dvss.n1835 9.3005
R12272 dvss.n1926 dvss.n1843 9.3005
R12273 dvss.n1925 dvss.n1844 9.3005
R12274 dvss.n1852 dvss.n1847 9.3005
R12275 dvss.n1915 dvss.n1848 9.3005
R12276 dvss.n1912 dvss.n698 9.3005
R12277 dvss.n3157 dvss.n3156 9.3005
R12278 dvss.n3161 dvss.n693 9.3005
R12279 dvss.n3183 dvss.n3182 9.3005
R12280 dvss.n3179 dvss.n694 9.3005
R12281 dvss.n3178 dvss.n3170 9.3005
R12282 dvss.n3177 dvss.n3176 9.3005
R12283 dvss.n3191 dvss.n684 9.3005
R12284 dvss.n683 dvss.n682 9.3005
R12285 dvss.n3198 dvss.n3197 9.3005
R12286 dvss.n3204 dvss.n678 9.3005
R12287 dvss.n3211 dvss.n3210 9.3005
R12288 dvss.n3217 dvss.n670 9.3005
R12289 dvss.n3226 dvss.n3225 9.3005
R12290 dvss.n3229 dvss.n3227 9.3005
R12291 dvss.n3228 dvss.n667 9.3005
R12292 dvss.n3241 dvss.n661 9.3005
R12293 dvss.n3247 dvss.n3246 9.3005
R12294 dvss.n3256 dvss.n3248 9.3005
R12295 dvss.n3255 dvss.n657 9.3005
R12296 dvss.n3274 dvss.n649 9.3005
R12297 dvss.n3271 dvss.n654 9.3005
R12298 dvss.n3270 dvss.n3269 9.3005
R12299 dvss.n3280 dvss.n640 9.3005
R12300 dvss.n3284 dvss.n3283 9.3005
R12301 dvss.n642 dvss.n634 9.3005
R12302 dvss.n3303 dvss.n3302 9.3005
R12303 dvss.n3299 dvss.n635 9.3005
R12304 dvss.n3298 dvss.n628 9.3005
R12305 dvss.n3310 dvss.n3309 9.3005
R12306 dvss.n3316 dvss.n623 9.3005
R12307 dvss.n3320 dvss.n3319 9.3005
R12308 dvss.n624 dvss.n618 9.3005
R12309 dvss.n3330 dvss.n3329 9.3005
R12310 dvss.n3342 dvss.n613 9.3005
R12311 dvss.n3346 dvss.n3345 9.3005
R12312 dvss.n3336 dvss.n606 9.3005
R12313 dvss.n3354 dvss.n3353 9.3005
R12314 dvss.n3357 dvss.n602 9.3005
R12315 dvss.n3363 dvss.n3362 9.3005
R12316 dvss.n3369 dvss.n597 9.3005
R12317 dvss.n3377 dvss.n3376 9.3005
R12318 dvss.n3391 dvss.n586 9.3005
R12319 dvss.n3388 dvss.n3386 9.3005
R12320 dvss.n3387 dvss.n580 9.3005
R12321 dvss.n3398 dvss.n3397 9.3005
R12322 dvss.n3401 dvss.n3399 9.3005
R12323 dvss.n3400 dvss.n575 9.3005
R12324 dvss.n3415 dvss.n568 9.3005
R12325 dvss.n3414 dvss.n569 9.3005
R12326 dvss.n3413 dvss.n3412 9.3005
R12327 dvss.n3423 dvss.n559 9.3005
R12328 dvss.n3430 dvss.n3429 9.3005
R12329 dvss.n3438 dvss.n3431 9.3005
R12330 dvss.n3433 dvss.n556 9.3005
R12331 dvss.n3448 dvss.n550 9.3005
R12332 dvss.n3449 dvss.n545 9.3005
R12333 dvss.n3462 dvss.n3461 9.3005
R12334 dvss.n3458 dvss.n546 9.3005
R12335 dvss.n3457 dvss.n541 9.3005
R12336 dvss.n3473 dvss.n535 9.3005
R12337 dvss.n3479 dvss.n3478 9.3005
R12338 dvss.n3488 dvss.n3480 9.3005
R12339 dvss.n3487 dvss.n531 9.3005
R12340 dvss.n3505 dvss.n523 9.3005
R12341 dvss.n3502 dvss.n528 9.3005
R12342 dvss.n3501 dvss.n3500 9.3005
R12343 dvss.n3511 dvss.n514 9.3005
R12344 dvss.n3621 dvss.n3620 9.3005
R12345 dvss.n3617 dvss.n515 9.3005
R12346 dvss.n3616 dvss.n3515 9.3005
R12347 dvss.n3615 dvss.n3516 9.3005
R12348 dvss.n3612 dvss.n3520 9.3005
R12349 dvss.n3611 dvss.n3521 9.3005
R12350 dvss.n3552 dvss.n3524 9.3005
R12351 dvss.n3607 dvss.n3525 9.3005
R12352 dvss.n3604 dvss.n3530 9.3005
R12353 dvss.n3549 dvss.n3548 9.3005
R12354 dvss.n3551 dvss.n3550 9.3005
R12355 dvss.n3598 dvss.n3536 9.3005
R12356 dvss.n3595 dvss.n3541 9.3005
R12357 dvss.n3594 dvss.n3585 9.3005
R12358 dvss.n3586 dvss.n374 9.3005
R12359 dvss.n3893 dvss.n3892 9.3005
R12360 dvss.n3889 dvss.n375 9.3005
R12361 dvss.n3888 dvss.n379 9.3005
R12362 dvss.n452 dvss.n382 9.3005
R12363 dvss.n454 dvss.n453 9.3005
R12364 dvss.n460 dvss.n441 9.3005
R12365 dvss.n462 dvss.n461 9.3005
R12366 dvss.n3876 dvss.n388 9.3005
R12367 dvss.n3873 dvss.n393 9.3005
R12368 dvss.n3872 dvss.n394 9.3005
R12369 dvss.n3871 dvss.n395 9.3005
R12370 dvss.n3868 dvss.n399 9.3005
R12371 dvss.n3867 dvss.n400 9.3005
R12372 dvss.n3819 dvss.n403 9.3005
R12373 dvss.n3863 dvss.n404 9.3005
R12374 dvss.n3860 dvss.n409 9.3005
R12375 dvss.n3827 dvss.n3826 9.3005
R12376 dvss.n3829 dvss.n3828 9.3005
R12377 dvss.n3854 dvss.n415 9.3005
R12378 dvss.n3851 dvss.n420 9.3005
R12379 dvss.n3850 dvss.n421 9.3005
R12380 dvss.n3842 dvss.n348 9.3005
R12381 dvss.n3935 dvss.n3934 9.3005
R12382 dvss.n3937 dvss.n342 9.3005
R12383 dvss.n3946 dvss.n3945 9.3005
R12384 dvss.n3956 dvss.n338 9.3005
R12385 dvss.n3953 dvss.n333 9.3005
R12386 dvss.n3964 dvss.n3963 9.3005
R12387 dvss.n3962 dvss.n323 9.3005
R12388 dvss.n3974 dvss.n3973 9.3005
R12389 dvss.n3977 dvss.n319 9.3005
R12390 dvss.n3979 dvss.n3978 9.3005
R12391 dvss.n3985 dvss.n313 9.3005
R12392 dvss.n1055 dvss.n914 9.3005
R12393 dvss.n1054 dvss.n915 9.3005
R12394 dvss.n1053 dvss.n916 9.3005
R12395 dvss.n971 dvss.n917 9.3005
R12396 dvss.n1048 dvss.n919 9.3005
R12397 dvss.n1047 dvss.n920 9.3005
R12398 dvss.n1046 dvss.n921 9.3005
R12399 dvss.n982 dvss.n922 9.3005
R12400 dvss.n1040 dvss.n924 9.3005
R12401 dvss.n1039 dvss.n925 9.3005
R12402 dvss.n1038 dvss.n926 9.3005
R12403 dvss.n1008 dvss.n927 9.3005
R12404 dvss.n1032 dvss.n929 9.3005
R12405 dvss.n1031 dvss.n930 9.3005
R12406 dvss.n1030 dvss.n1029 9.3005
R12407 dvss.n934 dvss.n932 9.3005
R12408 dvss.n947 dvss.n946 9.3005
R12409 dvss.n948 dvss.n903 9.3005
R12410 dvss.n1238 dvss.n1237 9.3005
R12411 dvss.n1236 dvss.n901 9.3005
R12412 dvss.n1244 dvss.n897 9.3005
R12413 dvss.n1251 dvss.n1250 9.3005
R12414 dvss.n1257 dvss.n891 9.3005
R12415 dvss.n1264 dvss.n1263 9.3005
R12416 dvss.n1272 dvss.n887 9.3005
R12417 dvss.n1277 dvss.n1276 9.3005
R12418 dvss.n1275 dvss.n882 9.3005
R12419 dvss.n1288 dvss.n1287 9.3005
R12420 dvss.n1293 dvss.n878 9.3005
R12421 dvss.n1304 dvss.n1303 9.3005
R12422 dvss.n1302 dvss.n869 9.3005
R12423 dvss.n1320 dvss.n1319 9.3005
R12424 dvss.n1318 dvss.n1317 9.3005
R12425 dvss.n1316 dvss.n861 9.3005
R12426 dvss.n1327 dvss.n1326 9.3005
R12427 dvss.n1487 dvss.n1486 9.3005
R12428 dvss.n1485 dvss.n1484 9.3005
R12429 dvss.n1483 dvss.n1329 9.3005
R12430 dvss.n1482 dvss.n1481 9.3005
R12431 dvss.n1480 dvss.n1479 9.3005
R12432 dvss.n1478 dvss.n1334 9.3005
R12433 dvss.n1341 dvss.n1339 9.3005
R12434 dvss.n1474 dvss.n1473 9.3005
R12435 dvss.n1472 dvss.n1471 9.3005
R12436 dvss.n1409 dvss.n1344 9.3005
R12437 dvss.n1410 dvss.n1352 9.3005
R12438 dvss.n1465 dvss.n1464 9.3005
R12439 dvss.n1463 dvss.n1462 9.3005
R12440 dvss.n1461 dvss.n1355 9.3005
R12441 dvss.n1361 dvss.n1358 9.3005
R12442 dvss.n1454 dvss.n1453 9.3005
R12443 dvss.n1452 dvss.n1451 9.3005
R12444 dvss.n1450 dvss.n1364 9.3005
R12445 dvss.n1374 dvss.n1372 9.3005
R12446 dvss.n1440 dvss.n1439 9.3005
R12447 dvss.n1438 dvss.n1437 9.3005
R12448 dvss.n1679 dvss.n804 9.3005
R12449 dvss.n1684 dvss.n1683 9.3005
R12450 dvss.n1704 dvss.n1703 9.3005
R12451 dvss.n1702 dvss.n1701 9.3005
R12452 dvss.n1700 dvss.n1691 9.3005
R12453 dvss.n1699 dvss.n794 9.3005
R12454 dvss.n1713 dvss.n1712 9.3005
R12455 dvss.n1711 dvss.n792 9.3005
R12456 dvss.n1719 dvss.n788 9.3005
R12457 dvss.n1726 dvss.n1725 9.3005
R12458 dvss.n1732 dvss.n782 9.3005
R12459 dvss.n1739 dvss.n1738 9.3005
R12460 dvss.n1747 dvss.n778 9.3005
R12461 dvss.n1752 dvss.n1751 9.3005
R12462 dvss.n1750 dvss.n773 9.3005
R12463 dvss.n1763 dvss.n1762 9.3005
R12464 dvss.n1768 dvss.n769 9.3005
R12465 dvss.n1779 dvss.n1778 9.3005
R12466 dvss.n1777 dvss.n760 9.3005
R12467 dvss.n1795 dvss.n1794 9.3005
R12468 dvss.n1793 dvss.n1792 9.3005
R12469 dvss.n1791 dvss.n752 9.3005
R12470 dvss.n1802 dvss.n1801 9.3005
R12471 dvss.n1962 dvss.n1961 9.3005
R12472 dvss.n1960 dvss.n1959 9.3005
R12473 dvss.n1958 dvss.n1804 9.3005
R12474 dvss.n1957 dvss.n1956 9.3005
R12475 dvss.n1955 dvss.n1954 9.3005
R12476 dvss.n1953 dvss.n1809 9.3005
R12477 dvss.n1816 dvss.n1814 9.3005
R12478 dvss.n1949 dvss.n1948 9.3005
R12479 dvss.n1947 dvss.n1946 9.3005
R12480 dvss.n1884 dvss.n1819 9.3005
R12481 dvss.n1885 dvss.n1827 9.3005
R12482 dvss.n1940 dvss.n1939 9.3005
R12483 dvss.n1938 dvss.n1937 9.3005
R12484 dvss.n1936 dvss.n1830 9.3005
R12485 dvss.n1836 dvss.n1833 9.3005
R12486 dvss.n1929 dvss.n1928 9.3005
R12487 dvss.n1927 dvss.n1926 9.3005
R12488 dvss.n1925 dvss.n1839 9.3005
R12489 dvss.n1849 dvss.n1847 9.3005
R12490 dvss.n1915 dvss.n1914 9.3005
R12491 dvss.n1913 dvss.n1912 9.3005
R12492 dvss.n3157 dvss.n695 9.3005
R12493 dvss.n3162 dvss.n3161 9.3005
R12494 dvss.n3182 dvss.n3181 9.3005
R12495 dvss.n3180 dvss.n3179 9.3005
R12496 dvss.n3178 dvss.n3169 9.3005
R12497 dvss.n3177 dvss.n685 9.3005
R12498 dvss.n3191 dvss.n3190 9.3005
R12499 dvss.n3189 dvss.n683 9.3005
R12500 dvss.n3197 dvss.n679 9.3005
R12501 dvss.n3204 dvss.n3203 9.3005
R12502 dvss.n3210 dvss.n673 9.3005
R12503 dvss.n3217 dvss.n3216 9.3005
R12504 dvss.n3225 dvss.n669 9.3005
R12505 dvss.n3230 dvss.n3229 9.3005
R12506 dvss.n3228 dvss.n664 9.3005
R12507 dvss.n3241 dvss.n3240 9.3005
R12508 dvss.n3246 dvss.n660 9.3005
R12509 dvss.n3257 dvss.n3256 9.3005
R12510 dvss.n3255 dvss.n651 9.3005
R12511 dvss.n3274 dvss.n3273 9.3005
R12512 dvss.n3272 dvss.n3271 9.3005
R12513 dvss.n3270 dvss.n643 9.3005
R12514 dvss.n3281 dvss.n3280 9.3005
R12515 dvss.n3283 dvss.n3282 9.3005
R12516 dvss.n642 dvss.n636 9.3005
R12517 dvss.n3302 dvss.n3301 9.3005
R12518 dvss.n3300 dvss.n3299 9.3005
R12519 dvss.n3298 dvss.n3297 9.3005
R12520 dvss.n3310 dvss.n626 9.3005
R12521 dvss.n3317 dvss.n3316 9.3005
R12522 dvss.n3319 dvss.n3318 9.3005
R12523 dvss.n624 dvss.n621 9.3005
R12524 dvss.n3330 dvss.n614 9.3005
R12525 dvss.n3343 dvss.n3342 9.3005
R12526 dvss.n3345 dvss.n3344 9.3005
R12527 dvss.n3336 dvss.n604 9.3005
R12528 dvss.n3355 dvss.n3354 9.3005
R12529 dvss.n3357 dvss.n3356 9.3005
R12530 dvss.n3362 dvss.n598 9.3005
R12531 dvss.n3369 dvss.n3368 9.3005
R12532 dvss.n3376 dvss.n588 9.3005
R12533 dvss.n3391 dvss.n3390 9.3005
R12534 dvss.n3389 dvss.n3388 9.3005
R12535 dvss.n3387 dvss.n591 9.3005
R12536 dvss.n3397 dvss.n578 9.3005
R12537 dvss.n3402 dvss.n3401 9.3005
R12538 dvss.n3400 dvss.n566 9.3005
R12539 dvss.n3416 dvss.n3415 9.3005
R12540 dvss.n3414 dvss.n567 9.3005
R12541 dvss.n3413 dvss.n561 9.3005
R12542 dvss.n3423 dvss.n3422 9.3005
R12543 dvss.n3429 dvss.n558 9.3005
R12544 dvss.n3439 dvss.n3438 9.3005
R12545 dvss.n3433 dvss.n551 9.3005
R12546 dvss.n3448 dvss.n3447 9.3005
R12547 dvss.n3449 dvss.n547 9.3005
R12548 dvss.n3461 dvss.n3460 9.3005
R12549 dvss.n3459 dvss.n3458 9.3005
R12550 dvss.n3457 dvss.n538 9.3005
R12551 dvss.n3473 dvss.n3472 9.3005
R12552 dvss.n3478 dvss.n534 9.3005
R12553 dvss.n3489 dvss.n3488 9.3005
R12554 dvss.n3487 dvss.n525 9.3005
R12555 dvss.n3505 dvss.n3504 9.3005
R12556 dvss.n3503 dvss.n3502 9.3005
R12557 dvss.n3501 dvss.n517 9.3005
R12558 dvss.n3512 dvss.n3511 9.3005
R12559 dvss.n3620 dvss.n3619 9.3005
R12560 dvss.n3618 dvss.n3617 9.3005
R12561 dvss.n3616 dvss.n3514 9.3005
R12562 dvss.n3615 dvss.n3614 9.3005
R12563 dvss.n3613 dvss.n3612 9.3005
R12564 dvss.n3611 dvss.n3519 9.3005
R12565 dvss.n3526 dvss.n3524 9.3005
R12566 dvss.n3607 dvss.n3606 9.3005
R12567 dvss.n3605 dvss.n3604 9.3005
R12568 dvss.n3549 dvss.n3529 9.3005
R12569 dvss.n3550 dvss.n3537 9.3005
R12570 dvss.n3598 dvss.n3597 9.3005
R12571 dvss.n3596 dvss.n3595 9.3005
R12572 dvss.n3594 dvss.n3540 9.3005
R12573 dvss.n3586 dvss.n376 9.3005
R12574 dvss.n3892 dvss.n3891 9.3005
R12575 dvss.n3890 dvss.n3889 9.3005
R12576 dvss.n3888 dvss.n378 9.3005
R12577 dvss.n448 dvss.n382 9.3005
R12578 dvss.n453 dvss.n442 9.3005
R12579 dvss.n460 dvss.n459 9.3005
R12580 dvss.n461 dvss.n389 9.3005
R12581 dvss.n3876 dvss.n3875 9.3005
R12582 dvss.n3874 dvss.n3873 9.3005
R12583 dvss.n3872 dvss.n392 9.3005
R12584 dvss.n3871 dvss.n3870 9.3005
R12585 dvss.n3869 dvss.n3868 9.3005
R12586 dvss.n3867 dvss.n398 9.3005
R12587 dvss.n405 dvss.n403 9.3005
R12588 dvss.n3863 dvss.n3862 9.3005
R12589 dvss.n3861 dvss.n3860 9.3005
R12590 dvss.n3827 dvss.n408 9.3005
R12591 dvss.n3828 dvss.n416 9.3005
R12592 dvss.n3854 dvss.n3853 9.3005
R12593 dvss.n3852 dvss.n3851 9.3005
R12594 dvss.n3850 dvss.n419 9.3005
R12595 dvss.n3842 dvss.n3841 9.3005
R12596 dvss.n3935 dvss.n347 9.3005
R12597 dvss.n3938 dvss.n3937 9.3005
R12598 dvss.n3946 dvss.n340 9.3005
R12599 dvss.n3956 dvss.n3955 9.3005
R12600 dvss.n3954 dvss.n3953 9.3005
R12601 dvss.n3963 dvss.n331 9.3005
R12602 dvss.n3962 dvss.n320 9.3005
R12603 dvss.n3975 dvss.n3974 9.3005
R12604 dvss.n3977 dvss.n3976 9.3005
R12605 dvss.n3978 dvss.n314 9.3005
R12606 dvss.n3985 dvss.n3984 9.3005
R12607 dvss.n2869 dvss.n2868 9.3005
R12608 dvss.n2870 dvss.n2869 9.3005
R12609 dvss.n2861 dvss.n2860 9.3005
R12610 dvss.n2862 dvss.n2861 9.3005
R12611 dvss.n2850 dvss.n2849 9.3005
R12612 dvss.n2851 dvss.n2850 9.3005
R12613 dvss.n2816 dvss.n2815 9.3005
R12614 dvss.n2817 dvss.n2816 9.3005
R12615 dvss.n2825 dvss.n2823 9.3005
R12616 dvss.n2826 dvss.n2825 9.3005
R12617 dvss.n2833 dvss.n2831 9.3005
R12618 dvss.n2834 dvss.n2833 9.3005
R12619 dvss.n2803 dvss.n2802 9.3005
R12620 dvss.n2804 dvss.n2803 9.3005
R12621 dvss.n2769 dvss.n2768 9.3005
R12622 dvss.n2770 dvss.n2769 9.3005
R12623 dvss.n2778 dvss.n2776 9.3005
R12624 dvss.n2779 dvss.n2778 9.3005
R12625 dvss.n2786 dvss.n2784 9.3005
R12626 dvss.n2787 dvss.n2786 9.3005
R12627 dvss.n2756 dvss.n2755 9.3005
R12628 dvss.n2757 dvss.n2756 9.3005
R12629 dvss.n2722 dvss.n2721 9.3005
R12630 dvss.n2723 dvss.n2722 9.3005
R12631 dvss.n2731 dvss.n2729 9.3005
R12632 dvss.n2732 dvss.n2731 9.3005
R12633 dvss.n2739 dvss.n2737 9.3005
R12634 dvss.n2740 dvss.n2739 9.3005
R12635 dvss.n2709 dvss.n2708 9.3005
R12636 dvss.n2710 dvss.n2709 9.3005
R12637 dvss.n2675 dvss.n2674 9.3005
R12638 dvss.n2676 dvss.n2675 9.3005
R12639 dvss.n2684 dvss.n2682 9.3005
R12640 dvss.n2685 dvss.n2684 9.3005
R12641 dvss.n2692 dvss.n2690 9.3005
R12642 dvss.n2693 dvss.n2692 9.3005
R12643 dvss.n2662 dvss.n2661 9.3005
R12644 dvss.n2663 dvss.n2662 9.3005
R12645 dvss.n2628 dvss.n2627 9.3005
R12646 dvss.n2629 dvss.n2628 9.3005
R12647 dvss.n2637 dvss.n2635 9.3005
R12648 dvss.n2638 dvss.n2637 9.3005
R12649 dvss.n2645 dvss.n2643 9.3005
R12650 dvss.n2646 dvss.n2645 9.3005
R12651 dvss.n2615 dvss.n2614 9.3005
R12652 dvss.n2616 dvss.n2615 9.3005
R12653 dvss.n2928 dvss.n2927 9.3005
R12654 dvss.n2929 dvss.n2928 9.3005
R12655 dvss.n2924 dvss.n2310 9.3005
R12656 dvss.n2924 dvss.n2923 9.3005
R12657 dvss.n2907 dvss.n2309 9.3005
R12658 dvss.n2905 dvss.n2309 9.3005
R12659 dvss.n2956 dvss.n2955 9.3005
R12660 dvss.n2955 dvss.n2952 9.3005
R12661 dvss.n2286 dvss.n2285 9.3005
R12662 dvss.n2286 dvss.n2216 9.3005
R12663 dvss.n2231 dvss.n2215 9.3005
R12664 dvss.n2229 dvss.n2215 9.3005
R12665 dvss.n2982 dvss.n2981 9.3005
R12666 dvss.n2981 dvss.n2980 9.3005
R12667 dvss.n2273 dvss.n2272 9.3005
R12668 dvss.n2274 dvss.n2273 9.3005
R12669 dvss.n4113 dvss.n4112 9.3005
R12670 dvss.n4113 dvss.n271 9.3005
R12671 dvss.n363 dvss.n270 9.3005
R12672 dvss.n365 dvss.n270 9.3005
R12673 dvss.n4118 dvss.n4117 9.3005
R12674 dvss.n4117 dvss.n4116 9.3005
R12675 dvss.n4100 dvss.n4099 9.3005
R12676 dvss.n4101 dvss.n4100 9.3005
R12677 dvss.n4066 dvss.n4065 9.3005
R12678 dvss.n4067 dvss.n4066 9.3005
R12679 dvss.n4075 dvss.n4073 9.3005
R12680 dvss.n4076 dvss.n4075 9.3005
R12681 dvss.n4083 dvss.n4081 9.3005
R12682 dvss.n4084 dvss.n4083 9.3005
R12683 dvss.n2886 dvss.n2392 9.3005
R12684 dvss.n2885 dvss.n2884 9.3005
R12685 dvss.n2883 dvss.n2882 9.3005
R12686 dvss.n2881 dvss.n2395 9.3005
R12687 dvss.n2880 dvss.n2879 9.3005
R12688 dvss.n2878 dvss.n2877 9.3005
R12689 dvss.n2876 dvss.n2400 9.3005
R12690 dvss.n2875 dvss.n2874 9.3005
R12691 dvss.n2873 dvss.n2872 9.3005
R12692 dvss.n2871 dvss.n2403 9.3005
R12693 dvss.n2867 dvss.n2866 9.3005
R12694 dvss.n2865 dvss.n2864 9.3005
R12695 dvss.n2863 dvss.n2411 9.3005
R12696 dvss.n2416 dvss.n2415 9.3005
R12697 dvss.n2859 dvss.n2858 9.3005
R12698 dvss.n2857 dvss.n2856 9.3005
R12699 dvss.n2855 dvss.n2854 9.3005
R12700 dvss.n2853 dvss.n2852 9.3005
R12701 dvss.n2426 dvss.n2423 9.3005
R12702 dvss.n2848 dvss.n2847 9.3005
R12703 dvss.n2846 dvss.n2845 9.3005
R12704 dvss.n2844 dvss.n2429 9.3005
R12705 dvss.n2843 dvss.n2842 9.3005
R12706 dvss.n2841 dvss.n2840 9.3005
R12707 dvss.n2839 dvss.n2434 9.3005
R12708 dvss.n2838 dvss.n2837 9.3005
R12709 dvss.n2836 dvss.n2835 9.3005
R12710 dvss.n2439 dvss.n2437 9.3005
R12711 dvss.n2830 dvss.n2829 9.3005
R12712 dvss.n2828 dvss.n2827 9.3005
R12713 dvss.n2445 dvss.n2444 9.3005
R12714 dvss.n2822 dvss.n2821 9.3005
R12715 dvss.n2820 dvss.n2819 9.3005
R12716 dvss.n2818 dvss.n2448 9.3005
R12717 dvss.n2814 dvss.n2813 9.3005
R12718 dvss.n2812 dvss.n2811 9.3005
R12719 dvss.n2810 dvss.n2453 9.3005
R12720 dvss.n2809 dvss.n2808 9.3005
R12721 dvss.n2807 dvss.n2806 9.3005
R12722 dvss.n2805 dvss.n2456 9.3005
R12723 dvss.n2462 dvss.n2459 9.3005
R12724 dvss.n2801 dvss.n2800 9.3005
R12725 dvss.n2799 dvss.n2798 9.3005
R12726 dvss.n2797 dvss.n2465 9.3005
R12727 dvss.n2796 dvss.n2795 9.3005
R12728 dvss.n2794 dvss.n2793 9.3005
R12729 dvss.n2792 dvss.n2470 9.3005
R12730 dvss.n2791 dvss.n2790 9.3005
R12731 dvss.n2789 dvss.n2788 9.3005
R12732 dvss.n2475 dvss.n2473 9.3005
R12733 dvss.n2783 dvss.n2782 9.3005
R12734 dvss.n2781 dvss.n2780 9.3005
R12735 dvss.n2481 dvss.n2480 9.3005
R12736 dvss.n2775 dvss.n2774 9.3005
R12737 dvss.n2773 dvss.n2772 9.3005
R12738 dvss.n2771 dvss.n2484 9.3005
R12739 dvss.n2767 dvss.n2766 9.3005
R12740 dvss.n2765 dvss.n2764 9.3005
R12741 dvss.n2763 dvss.n2489 9.3005
R12742 dvss.n2762 dvss.n2761 9.3005
R12743 dvss.n2760 dvss.n2759 9.3005
R12744 dvss.n2758 dvss.n2492 9.3005
R12745 dvss.n2498 dvss.n2495 9.3005
R12746 dvss.n2754 dvss.n2753 9.3005
R12747 dvss.n2752 dvss.n2751 9.3005
R12748 dvss.n2750 dvss.n2501 9.3005
R12749 dvss.n2749 dvss.n2748 9.3005
R12750 dvss.n2747 dvss.n2746 9.3005
R12751 dvss.n2745 dvss.n2506 9.3005
R12752 dvss.n2744 dvss.n2743 9.3005
R12753 dvss.n2742 dvss.n2741 9.3005
R12754 dvss.n2511 dvss.n2509 9.3005
R12755 dvss.n2736 dvss.n2735 9.3005
R12756 dvss.n2734 dvss.n2733 9.3005
R12757 dvss.n2517 dvss.n2516 9.3005
R12758 dvss.n2728 dvss.n2727 9.3005
R12759 dvss.n2726 dvss.n2725 9.3005
R12760 dvss.n2724 dvss.n2520 9.3005
R12761 dvss.n2720 dvss.n2719 9.3005
R12762 dvss.n2718 dvss.n2717 9.3005
R12763 dvss.n2716 dvss.n2525 9.3005
R12764 dvss.n2715 dvss.n2714 9.3005
R12765 dvss.n2713 dvss.n2712 9.3005
R12766 dvss.n2711 dvss.n2528 9.3005
R12767 dvss.n2534 dvss.n2531 9.3005
R12768 dvss.n2707 dvss.n2706 9.3005
R12769 dvss.n2705 dvss.n2704 9.3005
R12770 dvss.n2703 dvss.n2537 9.3005
R12771 dvss.n2702 dvss.n2701 9.3005
R12772 dvss.n2700 dvss.n2699 9.3005
R12773 dvss.n2698 dvss.n2542 9.3005
R12774 dvss.n2697 dvss.n2696 9.3005
R12775 dvss.n2695 dvss.n2694 9.3005
R12776 dvss.n2547 dvss.n2545 9.3005
R12777 dvss.n2689 dvss.n2688 9.3005
R12778 dvss.n2687 dvss.n2686 9.3005
R12779 dvss.n2553 dvss.n2552 9.3005
R12780 dvss.n2681 dvss.n2680 9.3005
R12781 dvss.n2679 dvss.n2678 9.3005
R12782 dvss.n2677 dvss.n2556 9.3005
R12783 dvss.n2673 dvss.n2672 9.3005
R12784 dvss.n2671 dvss.n2670 9.3005
R12785 dvss.n2669 dvss.n2561 9.3005
R12786 dvss.n2668 dvss.n2667 9.3005
R12787 dvss.n2666 dvss.n2665 9.3005
R12788 dvss.n2664 dvss.n2564 9.3005
R12789 dvss.n2570 dvss.n2567 9.3005
R12790 dvss.n2660 dvss.n2659 9.3005
R12791 dvss.n2658 dvss.n2657 9.3005
R12792 dvss.n2656 dvss.n2573 9.3005
R12793 dvss.n2655 dvss.n2654 9.3005
R12794 dvss.n2653 dvss.n2652 9.3005
R12795 dvss.n2651 dvss.n2578 9.3005
R12796 dvss.n2650 dvss.n2649 9.3005
R12797 dvss.n2648 dvss.n2647 9.3005
R12798 dvss.n2583 dvss.n2581 9.3005
R12799 dvss.n2642 dvss.n2641 9.3005
R12800 dvss.n2640 dvss.n2639 9.3005
R12801 dvss.n2589 dvss.n2588 9.3005
R12802 dvss.n2634 dvss.n2633 9.3005
R12803 dvss.n2632 dvss.n2631 9.3005
R12804 dvss.n2630 dvss.n2592 9.3005
R12805 dvss.n2626 dvss.n2625 9.3005
R12806 dvss.n2624 dvss.n2623 9.3005
R12807 dvss.n2622 dvss.n2597 9.3005
R12808 dvss.n2621 dvss.n2620 9.3005
R12809 dvss.n2619 dvss.n2618 9.3005
R12810 dvss.n2617 dvss.n2600 9.3005
R12811 dvss.n2606 dvss.n2603 9.3005
R12812 dvss.n2613 dvss.n2612 9.3005
R12813 dvss.n2611 dvss.n2610 9.3005
R12814 dvss.n2609 dvss.n2323 9.3005
R12815 dvss.n2893 dvss.n2892 9.3005
R12816 dvss.n2894 dvss.n2322 9.3005
R12817 dvss.n2897 dvss.n2896 9.3005
R12818 dvss.n2895 dvss.n2318 9.3005
R12819 dvss.n2904 dvss.n2903 9.3005
R12820 dvss.n2906 dvss.n2317 9.3005
R12821 dvss.n2910 dvss.n2909 9.3005
R12822 dvss.n2908 dvss.n2312 9.3005
R12823 dvss.n2922 dvss.n2921 9.3005
R12824 dvss.n2920 dvss.n2919 9.3005
R12825 dvss.n2918 dvss.n2307 9.3005
R12826 dvss.n2931 dvss.n2930 9.3005
R12827 dvss.n2926 dvss.n2304 9.3005
R12828 dvss.n2939 dvss.n2938 9.3005
R12829 dvss.n2940 dvss.n2303 9.3005
R12830 dvss.n2943 dvss.n2942 9.3005
R12831 dvss.n2941 dvss.n2299 9.3005
R12832 dvss.n2951 dvss.n2950 9.3005
R12833 dvss.n2298 dvss.n2297 9.3005
R12834 dvss.n2959 dvss.n2958 9.3005
R12835 dvss.n2957 dvss.n2294 9.3005
R12836 dvss.n2966 dvss.n2965 9.3005
R12837 dvss.n2967 dvss.n2293 9.3005
R12838 dvss.n2970 dvss.n2969 9.3005
R12839 dvss.n2968 dvss.n2289 9.3005
R12840 dvss.n2978 dvss.n2977 9.3005
R12841 dvss.n2979 dvss.n2212 9.3005
R12842 dvss.n2984 dvss.n2983 9.3005
R12843 dvss.n2223 dvss.n2213 9.3005
R12844 dvss.n2228 dvss.n2227 9.3005
R12845 dvss.n2230 dvss.n2221 9.3005
R12846 dvss.n2235 dvss.n2234 9.3005
R12847 dvss.n2233 dvss.n2222 9.3005
R12848 dvss.n2232 dvss.n2217 9.3005
R12849 dvss.n2284 dvss.n2283 9.3005
R12850 dvss.n2282 dvss.n2281 9.3005
R12851 dvss.n2280 dvss.n2243 9.3005
R12852 dvss.n2279 dvss.n2278 9.3005
R12853 dvss.n2277 dvss.n2276 9.3005
R12854 dvss.n2275 dvss.n2246 9.3005
R12855 dvss.n2271 dvss.n2270 9.3005
R12856 dvss.n259 dvss.n258 9.3005
R12857 dvss.n4132 dvss.n4131 9.3005
R12858 dvss.n4130 dvss.n4129 9.3005
R12859 dvss.n4128 dvss.n262 9.3005
R12860 dvss.n4127 dvss.n4126 9.3005
R12861 dvss.n4125 dvss.n4124 9.3005
R12862 dvss.n4123 dvss.n265 9.3005
R12863 dvss.n4122 dvss.n4121 9.3005
R12864 dvss.n4120 dvss.n4119 9.3005
R12865 dvss.n358 dvss.n268 9.3005
R12866 dvss.n367 dvss.n366 9.3005
R12867 dvss.n364 dvss.n357 9.3005
R12868 dvss.n362 dvss.n361 9.3005
R12869 dvss.n360 dvss.n351 9.3005
R12870 dvss.n359 dvss.n272 9.3005
R12871 dvss.n4111 dvss.n4110 9.3005
R12872 dvss.n4109 dvss.n4108 9.3005
R12873 dvss.n4107 dvss.n275 9.3005
R12874 dvss.n4106 dvss.n4105 9.3005
R12875 dvss.n4104 dvss.n4103 9.3005
R12876 dvss.n4102 dvss.n278 9.3005
R12877 dvss.n282 dvss.n281 9.3005
R12878 dvss.n4098 dvss.n4097 9.3005
R12879 dvss.n4096 dvss.n4095 9.3005
R12880 dvss.n4094 dvss.n285 9.3005
R12881 dvss.n4093 dvss.n4092 9.3005
R12882 dvss.n4091 dvss.n4090 9.3005
R12883 dvss.n4089 dvss.n288 9.3005
R12884 dvss.n4088 dvss.n4087 9.3005
R12885 dvss.n4086 dvss.n4085 9.3005
R12886 dvss.n293 dvss.n291 9.3005
R12887 dvss.n4080 dvss.n4079 9.3005
R12888 dvss.n4078 dvss.n4077 9.3005
R12889 dvss.n297 dvss.n296 9.3005
R12890 dvss.n4072 dvss.n4071 9.3005
R12891 dvss.n4070 dvss.n4069 9.3005
R12892 dvss.n4068 dvss.n300 9.3005
R12893 dvss.n4064 dvss.n4063 9.3005
R12894 dvss.n4062 dvss.n4061 9.3005
R12895 dvss.n4060 dvss.n303 9.3005
R12896 dvss.n4059 dvss.n4058 9.3005
R12897 dvss.n144 dvss.n143 9.3005
R12898 dvss.n147 dvss.n146 9.3005
R12899 dvss.n148 dvss.n100 9.3005
R12900 dvss.n150 dvss.n149 9.3005
R12901 dvss.n151 dvss.n98 9.3005
R12902 dvss.n118 dvss.n117 9.3005
R12903 dvss.n119 dvss.n111 9.3005
R12904 dvss.n121 dvss.n120 9.3005
R12905 dvss.n123 dvss.n109 9.3005
R12906 dvss.n127 dvss.n126 9.3005
R12907 dvss.n128 dvss.n108 9.3005
R12908 dvss.n130 dvss.n129 9.3005
R12909 dvss.n132 dvss.n106 9.3005
R12910 dvss.n136 dvss.n135 9.3005
R12911 dvss.n138 dvss.n137 9.3005
R12912 dvss.n140 dvss.n102 9.3005
R12913 dvss.n142 dvss.n141 9.3005
R12914 dvss.n254 dvss.n6 9.3005
R12915 dvss.n253 dvss.n252 9.3005
R12916 dvss.n251 dvss.n8 9.3005
R12917 dvss.n250 dvss.n249 9.3005
R12918 dvss.n247 dvss.n246 9.3005
R12919 dvss.n26 dvss.n25 9.3005
R12920 dvss.n27 dvss.n19 9.3005
R12921 dvss.n29 dvss.n28 9.3005
R12922 dvss.n31 dvss.n17 9.3005
R12923 dvss.n35 dvss.n34 9.3005
R12924 dvss.n36 dvss.n16 9.3005
R12925 dvss.n38 dvss.n37 9.3005
R12926 dvss.n40 dvss.n14 9.3005
R12927 dvss.n239 dvss.n238 9.3005
R12928 dvss.n241 dvss.n240 9.3005
R12929 dvss.n243 dvss.n10 9.3005
R12930 dvss.n245 dvss.n244 9.3005
R12931 dvss.n164 dvss.n163 9.3005
R12932 dvss.n162 dvss.n161 9.3005
R12933 dvss.n160 dvss.n159 9.3005
R12934 dvss.n158 dvss.n95 9.3005
R12935 dvss.n157 dvss.n156 9.3005
R12936 dvss.n74 dvss.n73 9.3005
R12937 dvss.n76 dvss.n68 9.3005
R12938 dvss.n80 dvss.n79 9.3005
R12939 dvss.n81 dvss.n67 9.3005
R12940 dvss.n83 dvss.n82 9.3005
R12941 dvss.n85 dvss.n65 9.3005
R12942 dvss.n89 dvss.n88 9.3005
R12943 dvss.n90 dvss.n62 9.3005
R12944 dvss.n172 dvss.n171 9.3005
R12945 dvss.n170 dvss.n169 9.3005
R12946 dvss.n167 dvss.n91 9.3005
R12947 dvss.n166 dvss.n165 9.3005
R12948 dvss.n228 dvss.n227 9.3005
R12949 dvss.n226 dvss.n225 9.3005
R12950 dvss.n224 dvss.n223 9.3005
R12951 dvss.n222 dvss.n217 9.3005
R12952 dvss.n221 dvss.n220 9.3005
R12953 dvss.n2 dvss.n0 9.3005
R12954 dvss.n4143 dvss.n4142 9.3005
R12955 dvss.n4140 dvss.n1 9.3005
R12956 dvss.n4139 dvss.n4138 9.3005
R12957 dvss.n4137 dvss.n4 9.3005
R12958 dvss.n195 dvss.n194 9.3005
R12959 dvss.n196 dvss.n188 9.3005
R12960 dvss.n198 dvss.n197 9.3005
R12961 dvss.n200 dvss.n186 9.3005
R12962 dvss.n204 dvss.n203 9.3005
R12963 dvss.n205 dvss.n185 9.3005
R12964 dvss.n207 dvss.n206 9.3005
R12965 dvss.n209 dvss.n183 9.3005
R12966 dvss.n213 dvss.n212 9.3005
R12967 dvss.n214 dvss.n180 9.3005
R12968 dvss.n231 dvss.n230 9.3005
R12969 dvss.n229 dvss.n182 9.3005
R12970 dvss.n1023 dvss.n1021 8.56999
R12971 dvss.n2414 dvss.n2412 8.56999
R12972 dvss.n3865 dvss.n402 8.54791
R12973 dvss.n3609 dvss.n3523 8.54791
R12974 dvss.n3427 dvss.n3426 8.54791
R12975 dvss.n3314 dvss.n3313 8.54791
R12976 dvss.n3195 dvss.n3194 8.54791
R12977 dvss.n1951 dvss.n1813 8.54791
R12978 dvss.n1717 dvss.n1716 8.54791
R12979 dvss.n1476 dvss.n1338 8.54791
R12980 dvss.n1242 dvss.n1241 8.54791
R12981 dvss.n4100 dvss.n280 8.54791
R12982 dvss.n2273 dvss.n2248 8.54791
R12983 dvss.n2955 dvss.n2954 8.54791
R12984 dvss.n2615 dvss.n2602 8.54791
R12985 dvss.n2662 dvss.n2566 8.54791
R12986 dvss.n2709 dvss.n2530 8.54791
R12987 dvss.n2756 dvss.n2494 8.54791
R12988 dvss.n2803 dvss.n2458 8.54791
R12989 dvss.n2850 dvss.n2425 8.54791
R12990 dvss.n1003 dvss 8.48432
R12991 dvss.n2404 dvss 8.48432
R12992 dvss.n402 dvss 8.43944
R12993 dvss.n3523 dvss 8.43944
R12994 dvss.n3426 dvss 8.43944
R12995 dvss.n3313 dvss 8.43944
R12996 dvss.n3194 dvss 8.43944
R12997 dvss.n1813 dvss 8.43944
R12998 dvss.n1716 dvss 8.43944
R12999 dvss.n1338 dvss 8.43944
R13000 dvss.n1241 dvss 8.43944
R13001 dvss.n280 dvss 8.43944
R13002 dvss.n2248 dvss 8.43944
R13003 dvss.n2954 dvss 8.43944
R13004 dvss.n2602 dvss 8.43944
R13005 dvss.n2566 dvss 8.43944
R13006 dvss.n2530 dvss 8.43944
R13007 dvss.n2494 dvss 8.43944
R13008 dvss.n2458 dvss 8.43944
R13009 dvss.n2425 dvss 8.43944
R13010 dvss.n125 dvss.n108 8.35606
R13011 dvss.n85 dvss.n84 8.35606
R13012 dvss.n33 dvss.n16 8.2416
R13013 dvss.n126 dvss.n125 8.0005
R13014 dvss.n84 dvss.n83 8.0005
R13015 dvss.n1095 dvss.t277 7.99565
R13016 dvss.n34 dvss.n33 7.89091
R13017 dvss.n202 dvss.n185 7.5205
R13018 dvss.n1024 dvss.n1023 7.37677
R13019 dvss.n2861 dvss.n2414 7.37677
R13020 dvss.n4037 dvss.n3991 7.3244
R13021 dvss.n4045 dvss.n4044 7.25358
R13022 dvss.n203 dvss.n202 7.2005
R13023 dvss.n233 dvss.n232 7.2005
R13024 dvss.n233 dvss.n180 7.0405
R13025 dvss.n3738 dvss 6.4005
R13026 dvss.n478 dvss 6.4005
R13027 dvss.n2126 dvss 6.4005
R13028 dvss.n2095 dvss 6.4005
R13029 dvss.n2064 dvss 6.4005
R13030 dvss.n714 dvss 6.4005
R13031 dvss.n1589 dvss 6.4005
R13032 dvss.n823 dvss 6.4005
R13033 dvss.n1158 dvss 6.4005
R13034 dvss.n3951 dvss 6.4005
R13035 dvss.n380 dvss 6.4005
R13036 dvss.n3482 dvss 6.4005
R13037 dvss.n3371 dvss 6.4005
R13038 dvss.n3250 dvss 6.4005
R13039 dvss.n1845 dvss 6.4005
R13040 dvss.n1772 dvss 6.4005
R13041 dvss.n1370 dvss 6.4005
R13042 dvss.n1297 dvss 6.4005
R13043 dvss.n114 dvss.n112 5.90523
R13044 dvss.n72 dvss.n71 5.90523
R13045 dvss.n22 dvss.n20 5.87299
R13046 dvss dvss.n154 5.68051
R13047 dvss.n191 dvss.n189 5.65757
R13048 dvss.n123 dvss.n122 5.51161
R13049 dvss.n78 dvss.n67 5.51161
R13050 dvss.n3766 dvss 5.45235
R13051 dvss.n3687 dvss 5.45235
R13052 dvss.n3009 dvss 5.45235
R13053 dvss.n3059 dvss 5.45235
R13054 dvss.n3109 dvss 5.45235
R13055 dvss.n2029 dvss 5.45235
R13056 dvss.n1631 dvss 5.45235
R13057 dvss.n1554 dvss 5.45235
R13058 dvss.n1157 dvss 5.45235
R13059 dvss.n3950 dvss 5.45235
R13060 dvss.n3886 dvss 5.45235
R13061 dvss.n3485 dvss 5.45235
R13062 dvss.n3374 dvss 5.45235
R13063 dvss.n3253 dvss 5.45235
R13064 dvss.n1923 dvss 5.45235
R13065 dvss.n1775 dvss 5.45235
R13066 dvss.n1448 dvss 5.45235
R13067 dvss.n1300 dvss 5.45235
R13068 dvss.n31 dvss.n30 5.43612
R13069 dvss.n131 dvss.n130 5.15606
R13070 dvss.n88 dvss.n87 5.15606
R13071 dvss.n39 dvss.n38 5.08543
R13072 dvss.n200 dvss.n199 4.9605
R13073 dvss dvss.n4134 4.88722
R13074 dvss.n257 dvss 4.88201
R13075 dvss.n154 dvss 4.8781
R13076 dvss.n4046 dvss.n4045 4.80519
R13077 dvss.n208 dvss.n207 4.6405
R13078 dvss.n4032 dvss.n4008 4.58109
R13079 dvss.n4038 dvss.n4037 4.25273
R13080 dvss.n3959 dvss.n3958 3.68864
R13081 dvss.n3882 dvss.n3879 3.68864
R13082 dvss.n3508 dvss.n3507 3.68864
R13083 dvss.n3394 dvss.n3393 3.68864
R13084 dvss.n3277 dvss.n3276 3.68864
R13085 dvss.n1919 dvss.n697 3.68864
R13086 dvss.n1798 dvss.n1797 3.68864
R13087 dvss.n1444 dvss.n806 3.68864
R13088 dvss.n1323 dvss.n1322 3.68864
R13089 dvss.n4075 dvss.n292 3.68864
R13090 dvss.n4114 dvss.n270 3.68864
R13091 dvss.n2287 dvss.n2215 3.68864
R13092 dvss.n2925 dvss.n2924 3.68864
R13093 dvss.n2637 dvss.n2582 3.68864
R13094 dvss.n2684 dvss.n2546 3.68864
R13095 dvss.n2731 dvss.n2510 3.68864
R13096 dvss.n2778 dvss.n2474 3.68864
R13097 dvss.n2825 dvss.n2438 3.68864
R13098 dvss.n1021 dvss 3.25474
R13099 dvss.n2412 dvss 3.25474
R13100 dvss.n4134 dvss.n4133 2.94679
R13101 dvss.n3986 dvss 2.94111
R13102 dvss.n354 dvss.n352 2.87444
R13103 dvss.n3766 dvss.n3765 2.84494
R13104 dvss.n3688 dvss.n3687 2.84494
R13105 dvss.n3009 dvss.n3008 2.84494
R13106 dvss.n3059 dvss.n3058 2.84494
R13107 dvss.n3109 dvss.n3108 2.84494
R13108 dvss.n2030 dvss.n2029 2.84494
R13109 dvss.n1631 dvss.n1630 2.84494
R13110 dvss.n1555 dvss.n1554 2.84494
R13111 dvss.n1157 dvss.n1156 2.84494
R13112 dvss.n3950 dvss.n3949 2.84494
R13113 dvss.n3886 dvss.n3885 2.84494
R13114 dvss.n3485 dvss.n3484 2.84494
R13115 dvss.n3374 dvss.n3373 2.84494
R13116 dvss.n3253 dvss.n3252 2.84494
R13117 dvss.n1923 dvss.n1922 2.84494
R13118 dvss.n1775 dvss.n1774 2.84494
R13119 dvss.n1448 dvss.n1447 2.84494
R13120 dvss.n1300 dvss.n1299 2.84494
R13121 dvss.t266 dvss.t200 2.67324
R13122 dvss.n116 dvss.n111 2.66717
R13123 dvss.n76 dvss.n75 2.66717
R13124 dvss.n24 dvss.n19 2.63064
R13125 dvss.n3765 dvss 2.60791
R13126 dvss.n3688 dvss 2.60791
R13127 dvss.n3008 dvss 2.60791
R13128 dvss.n3058 dvss 2.60791
R13129 dvss.n3108 dvss 2.60791
R13130 dvss.n2030 dvss 2.60791
R13131 dvss.n1630 dvss 2.60791
R13132 dvss.n1555 dvss 2.60791
R13133 dvss.n1156 dvss 2.60791
R13134 dvss.n3949 dvss 2.60791
R13135 dvss.n3885 dvss 2.60791
R13136 dvss.n3484 dvss 2.60791
R13137 dvss.n3373 dvss 2.60791
R13138 dvss.n3252 dvss 2.60791
R13139 dvss.n1922 dvss 2.60791
R13140 dvss.n1774 dvss 2.60791
R13141 dvss.n1447 dvss 2.60791
R13142 dvss.n1299 dvss 2.60791
R13143 dvss.n1087 dvss 2.49542
R13144 dvss.n1075 dvss 2.49542
R13145 dvss.n1000 dvss 2.49542
R13146 dvss.n985 dvss 2.49542
R13147 dvss.n50 dvss.n5 2.43615
R13148 dvss.n4023 dvss.n4022 2.42979
R13149 dvss.n193 dvss.n188 2.4005
R13150 dvss.n135 dvss.n105 2.31161
R13151 dvss.n144 dvss.n101 2.31161
R13152 dvss.n172 dvss.n64 2.31161
R13153 dvss.n163 dvss.n93 2.31161
R13154 dvss.n238 dvss.n13 2.27995
R13155 dvss.n247 dvss.n9 2.27995
R13156 dvss.n48 dvss.n46 2.17238
R13157 dvss.n212 dvss.n211 2.0805
R13158 dvss.n227 dvss.n215 2.0805
R13159 dvss.n3775 dvss 1.84457
R13160 dvss dvss.n3774 1.84457
R13161 dvss.n3774 dvss 1.84457
R13162 dvss.n3673 dvss 1.84457
R13163 dvss dvss.n3672 1.84457
R13164 dvss.n3672 dvss 1.84457
R13165 dvss.n3018 dvss 1.84457
R13166 dvss dvss.n3017 1.84457
R13167 dvss.n3017 dvss 1.84457
R13168 dvss.n3068 dvss 1.84457
R13169 dvss dvss.n3067 1.84457
R13170 dvss.n3067 dvss 1.84457
R13171 dvss.n3118 dvss 1.84457
R13172 dvss dvss.n3117 1.84457
R13173 dvss.n3117 dvss 1.84457
R13174 dvss.n2015 dvss 1.84457
R13175 dvss dvss.n2014 1.84457
R13176 dvss.n2014 dvss 1.84457
R13177 dvss.n1640 dvss 1.84457
R13178 dvss dvss.n1639 1.84457
R13179 dvss.n1639 dvss 1.84457
R13180 dvss.n1540 dvss 1.84457
R13181 dvss dvss.n1539 1.84457
R13182 dvss.n1539 dvss 1.84457
R13183 dvss.n1143 dvss 1.84457
R13184 dvss dvss.n1140 1.84457
R13185 dvss.n1140 dvss 1.84457
R13186 dvss.n3848 dvss 1.84457
R13187 dvss dvss.n3847 1.84457
R13188 dvss.n3847 dvss 1.84457
R13189 dvss.n3592 dvss 1.84457
R13190 dvss dvss.n3591 1.84457
R13191 dvss.n3591 dvss 1.84457
R13192 dvss.n3475 dvss 1.84457
R13193 dvss.n3454 dvss 1.84457
R13194 dvss.n3454 dvss 1.84457
R13195 dvss.n3359 dvss 1.84457
R13196 dvss.n3335 dvss 1.84457
R13197 dvss.n3335 dvss 1.84457
R13198 dvss.n3243 dvss 1.84457
R13199 dvss.n3222 dvss 1.84457
R13200 dvss.n3222 dvss 1.84457
R13201 dvss.n1934 dvss 1.84457
R13202 dvss dvss.n1933 1.84457
R13203 dvss.n1933 dvss 1.84457
R13204 dvss.n1765 dvss 1.84457
R13205 dvss.n1744 dvss 1.84457
R13206 dvss.n1744 dvss 1.84457
R13207 dvss.n1459 dvss 1.84457
R13208 dvss dvss.n1458 1.84457
R13209 dvss.n1458 dvss 1.84457
R13210 dvss.n1290 dvss 1.84457
R13211 dvss.n1269 dvss 1.84457
R13212 dvss.n1269 dvss 1.84457
R13213 dvss.n4028 dvss.n4014 1.81727
R13214 dvss.n4015 dvss.n4008 1.81727
R13215 dvss.n4046 dvss.n3986 1.5923
R13216 dvss.n237 dvss.n40 1.57858
R13217 dvss.n146 dvss.n145 1.42272
R13218 dvss.n162 dvss.n94 1.42272
R13219 dvss.n249 dvss.n248 1.40324
R13220 dvss.n3997 dvss.n3988 1.35909
R13221 dvss.n3792 dvss.n3791 1.34003
R13222 dvss.n3784 dvss.n3783 1.34003
R13223 dvss.n3783 dvss.n3782 1.34003
R13224 dvss.n3656 dvss.n495 1.34003
R13225 dvss.n3658 dvss.n486 1.34003
R13226 dvss.n3671 dvss.n486 1.34003
R13227 dvss.n3035 dvss.n3034 1.34003
R13228 dvss.n3027 dvss.n3026 1.34003
R13229 dvss.n3026 dvss.n3025 1.34003
R13230 dvss.n3085 dvss.n3084 1.34003
R13231 dvss.n3077 dvss.n3076 1.34003
R13232 dvss.n3076 dvss.n3075 1.34003
R13233 dvss.n3135 dvss.n3134 1.34003
R13234 dvss.n3127 dvss.n3126 1.34003
R13235 dvss.n3126 dvss.n3125 1.34003
R13236 dvss.n1998 dvss.n731 1.34003
R13237 dvss.n2000 dvss.n722 1.34003
R13238 dvss.n2013 dvss.n722 1.34003
R13239 dvss.n1657 dvss.n1656 1.34003
R13240 dvss.n1649 dvss.n1648 1.34003
R13241 dvss.n1648 dvss.n1647 1.34003
R13242 dvss.n1523 dvss.n840 1.34003
R13243 dvss.n1525 dvss.n831 1.34003
R13244 dvss.n1538 dvss.n831 1.34003
R13245 dvss.n1131 dvss.n1129 1.34003
R13246 dvss.n1137 dvss.n1135 1.34003
R13247 dvss.n1139 dvss.n1137 1.34003
R13248 dvss.n3858 dvss.n412 1.34003
R13249 dvss.n3856 dvss.n414 1.34003
R13250 dvss.n3846 dvss.n414 1.34003
R13251 dvss.n3602 dvss.n3533 1.34003
R13252 dvss.n3600 dvss.n3535 1.34003
R13253 dvss.n3590 dvss.n3535 1.34003
R13254 dvss.n3436 dvss.n3435 1.34003
R13255 dvss.n3453 dvss.n3451 1.34003
R13256 dvss.n3455 dvss.n3453 1.34003
R13257 dvss.n3332 dvss.n617 1.34003
R13258 dvss.n3340 dvss.n3339 1.34003
R13259 dvss.n3339 dvss.n3338 1.34003
R13260 dvss.n3208 dvss.n3207 1.34003
R13261 dvss.n3221 dvss.n3219 1.34003
R13262 dvss.n3223 dvss.n3221 1.34003
R13263 dvss.n1944 dvss.n1823 1.34003
R13264 dvss.n1942 dvss.n1825 1.34003
R13265 dvss.n1932 dvss.n1825 1.34003
R13266 dvss.n1730 dvss.n1729 1.34003
R13267 dvss.n1743 dvss.n1741 1.34003
R13268 dvss.n1745 dvss.n1743 1.34003
R13269 dvss.n1469 dvss.n1348 1.34003
R13270 dvss.n1467 dvss.n1350 1.34003
R13271 dvss.n1457 dvss.n1350 1.34003
R13272 dvss.n1255 dvss.n1254 1.34003
R13273 dvss.n1268 dvss.n1266 1.34003
R13274 dvss.n1270 dvss.n1268 1.34003
R13275 dvss.n226 dvss.n216 1.2805
R13276 dvss.n4142 dvss.n4141 1.2805
R13277 dvss dvss.n4046 1.23235
R13278 dvss.n257 dvss.n5 1.16554
R13279 dvss.n195 dvss.n189 1.12105
R13280 dvss.n4038 dvss.n3988 1.09648
R13281 dvss.n50 dvss.n49 1.09487
R13282 dvss.n26 dvss.n20 1.05227
R13283 dvss.n118 dvss.n112 1.04213
R13284 dvss.n73 dvss.n72 1.04213
R13285 dvss.n219 dvss.n2 0.9605
R13286 dvss.n154 dvss.n5 0.934094
R13287 dvss.n51 dvss.n50 0.886661
R13288 dvss.n3791 dvss 0.856314
R13289 dvss.n3784 dvss.n3712 0.856314
R13290 dvss.n3782 dvss 0.856314
R13291 dvss dvss.n3656 0.856314
R13292 dvss.n3658 dvss.n3657 0.856314
R13293 dvss dvss.n3671 0.856314
R13294 dvss.n3034 dvss 0.856314
R13295 dvss.n3027 dvss.n2116 0.856314
R13296 dvss.n3025 dvss 0.856314
R13297 dvss.n3084 dvss 0.856314
R13298 dvss.n3077 dvss.n2085 0.856314
R13299 dvss.n3075 dvss 0.856314
R13300 dvss.n3134 dvss 0.856314
R13301 dvss.n3127 dvss.n2054 0.856314
R13302 dvss.n3125 dvss 0.856314
R13303 dvss dvss.n1998 0.856314
R13304 dvss.n2000 dvss.n1999 0.856314
R13305 dvss dvss.n2013 0.856314
R13306 dvss.n1656 dvss 0.856314
R13307 dvss.n1649 dvss.n1579 0.856314
R13308 dvss.n1647 dvss 0.856314
R13309 dvss dvss.n1523 0.856314
R13310 dvss.n1525 dvss.n1524 0.856314
R13311 dvss dvss.n1538 0.856314
R13312 dvss dvss.n1131 0.856314
R13313 dvss.n1135 dvss.n1132 0.856314
R13314 dvss dvss.n1139 0.856314
R13315 dvss.n3858 dvss 0.856314
R13316 dvss.n3857 dvss.n3856 0.856314
R13317 dvss dvss.n3846 0.856314
R13318 dvss.n3602 dvss 0.856314
R13319 dvss.n3601 dvss.n3600 0.856314
R13320 dvss dvss.n3590 0.856314
R13321 dvss.n3435 dvss 0.856314
R13322 dvss.n3451 dvss.n549 0.856314
R13323 dvss.n3455 dvss 0.856314
R13324 dvss dvss.n3332 0.856314
R13325 dvss.n3340 dvss.n3333 0.856314
R13326 dvss.n3338 dvss 0.856314
R13327 dvss.n3208 dvss 0.856314
R13328 dvss.n3219 dvss.n672 0.856314
R13329 dvss.n3223 dvss 0.856314
R13330 dvss.n1944 dvss 0.856314
R13331 dvss.n1943 dvss.n1942 0.856314
R13332 dvss dvss.n1932 0.856314
R13333 dvss.n1730 dvss 0.856314
R13334 dvss.n1741 dvss.n781 0.856314
R13335 dvss.n1745 dvss 0.856314
R13336 dvss.n1469 dvss 0.856314
R13337 dvss.n1468 dvss.n1467 0.856314
R13338 dvss dvss.n1457 0.856314
R13339 dvss.n1255 dvss 0.856314
R13340 dvss.n1266 dvss.n890 0.856314
R13341 dvss.n1270 dvss 0.856314
R13342 dvss.n49 dvss.n44 0.7755
R13343 dvss.n57 dvss.n53 0.7755
R13344 dvss.n134 dvss.n132 0.711611
R13345 dvss.n173 dvss.n62 0.711611
R13346 dvss.n52 dvss.n51 0.705857
R13347 dvss.n4042 dvss.t652 0.627052
R13348 dvss.n4040 dvss.t223 0.627052
R13349 dvss.n4016 dvss.t480 0.627052
R13350 dvss.n4041 dvss.n4040 0.5805
R13351 dvss.n4043 dvss.n4042 0.5805
R13352 dvss.n4020 dvss.n4019 0.5805
R13353 dvss.n4019 dvss.n4018 0.5805
R13354 dvss.n4018 dvss.n4017 0.5805
R13355 dvss.n4017 dvss.n4016 0.5805
R13356 dvss.n4026 dvss.n3987 0.54848
R13357 dvss.n3986 dvss 0.543548
R13358 dvss.n140 dvss.n139 0.533833
R13359 dvss.n168 dvss.n167 0.533833
R13360 dvss.n53 dvss.n46 0.529518
R13361 dvss.n243 dvss.n242 0.526527
R13362 dvss.n4134 dvss 0.506359
R13363 dvss.n232 dvss.n231 0.4805
R13364 dvss.n4001 dvss.n4000 0.427268
R13365 dvss.n4004 dvss.n3991 0.312562
R13366 dvss.n3999 dvss.n3998 0.299742
R13367 dvss.n4044 dvss.n4041 0.279444
R13368 dvss.n4044 dvss.n4043 0.268206
R13369 dvss.n4005 dvss.n4004 0.254288
R13370 dvss.n49 dvss.n48 0.2505
R13371 dvss dvss.n257 0.187023
R13372 dvss.n4029 dvss.n4023 0.179346
R13373 dvss.n4027 dvss.n4026 0.179346
R13374 dvss.n4037 dvss.n4036 0.179346
R13375 dvss.n4006 dvss.n4005 0.179346
R13376 dvss.n53 dvss.n52 0.176839
R13377 dvss.n3991 dvss.n3990 0.174082
R13378 dvss.n4005 dvss.n4001 0.145702
R13379 dvss.n4026 dvss.n4025 0.129288
R13380 dvss.n119 dvss.n118 0.120292
R13381 dvss.n120 dvss.n119 0.120292
R13382 dvss.n120 dvss.n109 0.120292
R13383 dvss.n127 dvss.n109 0.120292
R13384 dvss.n128 dvss.n127 0.120292
R13385 dvss.n129 dvss.n128 0.120292
R13386 dvss.n129 dvss.n106 0.120292
R13387 dvss.n136 dvss.n106 0.120292
R13388 dvss.n137 dvss.n136 0.120292
R13389 dvss.n137 dvss.n102 0.120292
R13390 dvss.n142 dvss.n102 0.120292
R13391 dvss.n143 dvss.n142 0.120292
R13392 dvss.n148 dvss.n147 0.120292
R13393 dvss.n149 dvss.n148 0.120292
R13394 dvss.n149 dvss.n98 0.120292
R13395 dvss.n153 dvss.n98 0.120292
R13396 dvss.n27 dvss.n26 0.120292
R13397 dvss.n28 dvss.n27 0.120292
R13398 dvss.n28 dvss.n17 0.120292
R13399 dvss.n35 dvss.n17 0.120292
R13400 dvss.n36 dvss.n35 0.120292
R13401 dvss.n37 dvss.n36 0.120292
R13402 dvss.n37 dvss.n14 0.120292
R13403 dvss.n239 dvss.n14 0.120292
R13404 dvss.n240 dvss.n239 0.120292
R13405 dvss.n240 dvss.n10 0.120292
R13406 dvss.n245 dvss.n10 0.120292
R13407 dvss.n246 dvss.n245 0.120292
R13408 dvss.n251 dvss.n250 0.120292
R13409 dvss.n252 dvss.n251 0.120292
R13410 dvss.n252 dvss.n6 0.120292
R13411 dvss.n256 dvss.n6 0.120292
R13412 dvss.n73 dvss.n68 0.120292
R13413 dvss.n80 dvss.n68 0.120292
R13414 dvss.n81 dvss.n80 0.120292
R13415 dvss.n82 dvss.n81 0.120292
R13416 dvss.n82 dvss.n65 0.120292
R13417 dvss.n89 dvss.n65 0.120292
R13418 dvss.n90 dvss.n89 0.120292
R13419 dvss.n171 dvss.n90 0.120292
R13420 dvss.n171 dvss.n170 0.120292
R13421 dvss.n170 dvss.n91 0.120292
R13422 dvss.n165 dvss.n91 0.120292
R13423 dvss.n165 dvss.n164 0.120292
R13424 dvss.n161 dvss.n160 0.120292
R13425 dvss.n160 dvss.n95 0.120292
R13426 dvss.n156 dvss.n95 0.120292
R13427 dvss.n156 dvss.n155 0.120292
R13428 dvss.n196 dvss.n195 0.120292
R13429 dvss.n197 dvss.n196 0.120292
R13430 dvss.n197 dvss.n186 0.120292
R13431 dvss.n204 dvss.n186 0.120292
R13432 dvss.n205 dvss.n204 0.120292
R13433 dvss.n206 dvss.n205 0.120292
R13434 dvss.n206 dvss.n183 0.120292
R13435 dvss.n213 dvss.n183 0.120292
R13436 dvss.n214 dvss.n213 0.120292
R13437 dvss.n230 dvss.n214 0.120292
R13438 dvss.n230 dvss.n229 0.120292
R13439 dvss.n229 dvss.n228 0.120292
R13440 dvss.n225 dvss.n224 0.120292
R13441 dvss.n224 dvss.n217 0.120292
R13442 dvss.n220 dvss.n217 0.120292
R13443 dvss.n220 dvss.n0 0.120292
R13444 dvss.n4143 dvss.n1 0.120292
R13445 dvss.n4138 dvss.n1 0.120292
R13446 dvss.n4138 dvss.n4137 0.120292
R13447 dvss.n4137 dvss.n4136 0.120292
R13448 dvss.n4004 dvss.n4003 0.101043
R13449 dvss.n3998 dvss.n3997 0.100247
R13450 dvss.n4000 dvss.n3999 0.0989849
R13451 dvss.n4025 dvss.n3988 0.0888838
R13452 dvss.n4039 dvss.n3987 0.0808571
R13453 dvss dvss.n2886 0.067223
R13454 dvss dvss.n2885 0.067223
R13455 dvss.n2882 dvss 0.067223
R13456 dvss dvss.n2881 0.067223
R13457 dvss dvss.n2880 0.067223
R13458 dvss.n2877 dvss 0.067223
R13459 dvss dvss.n2876 0.067223
R13460 dvss dvss.n2875 0.067223
R13461 dvss.n2872 dvss 0.067223
R13462 dvss dvss.n2871 0.067223
R13463 dvss.n2864 dvss 0.067223
R13464 dvss dvss.n2863 0.067223
R13465 dvss.n2856 dvss 0.067223
R13466 dvss.n2852 dvss 0.067223
R13467 dvss.n2845 dvss 0.067223
R13468 dvss dvss.n2844 0.067223
R13469 dvss dvss.n2843 0.067223
R13470 dvss.n2840 dvss 0.067223
R13471 dvss dvss.n2839 0.067223
R13472 dvss dvss.n2838 0.067223
R13473 dvss.n2835 dvss 0.067223
R13474 dvss.n2827 dvss 0.067223
R13475 dvss.n2819 dvss 0.067223
R13476 dvss dvss.n2818 0.067223
R13477 dvss.n2811 dvss 0.067223
R13478 dvss dvss.n2810 0.067223
R13479 dvss dvss.n2809 0.067223
R13480 dvss dvss.n2805 0.067223
R13481 dvss.n2798 dvss 0.067223
R13482 dvss dvss.n2797 0.067223
R13483 dvss dvss.n2796 0.067223
R13484 dvss.n2793 dvss 0.067223
R13485 dvss dvss.n2792 0.067223
R13486 dvss dvss.n2791 0.067223
R13487 dvss.n2788 dvss 0.067223
R13488 dvss.n2780 dvss 0.067223
R13489 dvss.n2772 dvss 0.067223
R13490 dvss dvss.n2771 0.067223
R13491 dvss.n2764 dvss 0.067223
R13492 dvss dvss.n2763 0.067223
R13493 dvss dvss.n2762 0.067223
R13494 dvss dvss.n2758 0.067223
R13495 dvss.n2751 dvss 0.067223
R13496 dvss dvss.n2750 0.067223
R13497 dvss dvss.n2749 0.067223
R13498 dvss.n2746 dvss 0.067223
R13499 dvss dvss.n2745 0.067223
R13500 dvss dvss.n2744 0.067223
R13501 dvss.n2741 dvss 0.067223
R13502 dvss.n2733 dvss 0.067223
R13503 dvss.n2725 dvss 0.067223
R13504 dvss dvss.n2724 0.067223
R13505 dvss.n2717 dvss 0.067223
R13506 dvss dvss.n2716 0.067223
R13507 dvss dvss.n2715 0.067223
R13508 dvss dvss.n2711 0.067223
R13509 dvss.n2704 dvss 0.067223
R13510 dvss dvss.n2703 0.067223
R13511 dvss dvss.n2702 0.067223
R13512 dvss.n2699 dvss 0.067223
R13513 dvss dvss.n2698 0.067223
R13514 dvss dvss.n2697 0.067223
R13515 dvss.n2694 dvss 0.067223
R13516 dvss.n2686 dvss 0.067223
R13517 dvss.n2678 dvss 0.067223
R13518 dvss dvss.n2677 0.067223
R13519 dvss.n2670 dvss 0.067223
R13520 dvss dvss.n2669 0.067223
R13521 dvss dvss.n2668 0.067223
R13522 dvss dvss.n2664 0.067223
R13523 dvss.n2657 dvss 0.067223
R13524 dvss dvss.n2656 0.067223
R13525 dvss dvss.n2655 0.067223
R13526 dvss.n2652 dvss 0.067223
R13527 dvss dvss.n2651 0.067223
R13528 dvss dvss.n2650 0.067223
R13529 dvss.n2647 dvss 0.067223
R13530 dvss.n2639 dvss 0.067223
R13531 dvss.n2631 dvss 0.067223
R13532 dvss dvss.n2630 0.067223
R13533 dvss.n2623 dvss 0.067223
R13534 dvss dvss.n2622 0.067223
R13535 dvss dvss.n2621 0.067223
R13536 dvss dvss.n2617 0.067223
R13537 dvss.n2610 dvss 0.067223
R13538 dvss dvss.n2609 0.067223
R13539 dvss.n2893 dvss 0.067223
R13540 dvss.n2894 dvss 0.067223
R13541 dvss.n2896 dvss 0.067223
R13542 dvss dvss.n2895 0.067223
R13543 dvss.n2904 dvss 0.067223
R13544 dvss dvss.n2908 0.067223
R13545 dvss dvss.n2918 0.067223
R13546 dvss.n2930 dvss 0.067223
R13547 dvss.n2939 dvss 0.067223
R13548 dvss.n2940 dvss 0.067223
R13549 dvss.n2942 dvss 0.067223
R13550 dvss.n2951 dvss 0.067223
R13551 dvss dvss.n2957 0.067223
R13552 dvss.n2966 dvss 0.067223
R13553 dvss.n2967 dvss 0.067223
R13554 dvss.n2969 dvss 0.067223
R13555 dvss dvss.n2968 0.067223
R13556 dvss.n2978 dvss 0.067223
R13557 dvss.n2979 dvss 0.067223
R13558 dvss.n2228 dvss 0.067223
R13559 dvss dvss.n2233 0.067223
R13560 dvss dvss.n2232 0.067223
R13561 dvss.n2281 dvss 0.067223
R13562 dvss dvss.n2280 0.067223
R13563 dvss dvss.n2279 0.067223
R13564 dvss dvss.n2275 0.067223
R13565 dvss dvss.n4132 0.067223
R13566 dvss.n4129 dvss 0.067223
R13567 dvss dvss.n4128 0.067223
R13568 dvss dvss.n4127 0.067223
R13569 dvss.n4124 dvss 0.067223
R13570 dvss dvss.n4123 0.067223
R13571 dvss dvss.n4122 0.067223
R13572 dvss.n366 dvss 0.067223
R13573 dvss dvss.n360 0.067223
R13574 dvss dvss.n359 0.067223
R13575 dvss.n4108 dvss 0.067223
R13576 dvss dvss.n4107 0.067223
R13577 dvss dvss.n4106 0.067223
R13578 dvss dvss.n4102 0.067223
R13579 dvss.n4095 dvss 0.067223
R13580 dvss dvss.n4094 0.067223
R13581 dvss dvss.n4093 0.067223
R13582 dvss.n4090 dvss 0.067223
R13583 dvss dvss.n4089 0.067223
R13584 dvss dvss.n4088 0.067223
R13585 dvss.n4085 dvss 0.067223
R13586 dvss.n4077 dvss 0.067223
R13587 dvss.n4069 dvss 0.067223
R13588 dvss dvss.n4068 0.067223
R13589 dvss.n4061 dvss 0.067223
R13590 dvss dvss.n4060 0.067223
R13591 dvss dvss.n4059 0.067223
R13592 dvss dvss.n2826 0.0638446
R13593 dvss dvss.n2779 0.0638446
R13594 dvss dvss.n2732 0.0638446
R13595 dvss dvss.n2685 0.0638446
R13596 dvss dvss.n2638 0.0638446
R13597 dvss.n2923 dvss 0.0638446
R13598 dvss.n2229 dvss 0.0638446
R13599 dvss dvss.n365 0.0638446
R13600 dvss dvss.n4076 0.0638446
R13601 dvss dvss.n2848 0.0613108
R13602 dvss dvss.n2801 0.0613108
R13603 dvss dvss.n2754 0.0613108
R13604 dvss dvss.n2707 0.0613108
R13605 dvss dvss.n2660 0.0613108
R13606 dvss dvss.n2613 0.0613108
R13607 dvss.n2958 dvss 0.0613108
R13608 dvss dvss.n258 0.0613108
R13609 dvss dvss.n4098 0.0613108
R13610 dvss.n147 dvss 0.0603958
R13611 dvss.n250 dvss 0.0603958
R13612 dvss.n161 dvss 0.0603958
R13613 dvss.n225 dvss 0.0603958
R13614 dvss dvss.n4143 0.0603958
R13615 dvss.n4043 dvss.t222 0.047052
R13616 dvss.n4042 dvss.t654 0.047052
R13617 dvss.n4040 dvss.t655 0.047052
R13618 dvss.n4041 dvss.t653 0.047052
R13619 dvss.n4016 dvss.t479 0.047052
R13620 dvss.n4017 dvss.t488 0.047052
R13621 dvss.n4018 dvss.t483 0.047052
R13622 dvss.n4019 dvss.t485 0.047052
R13623 dvss.n4020 dvss.t484 0.047052
R13624 dvss.n2868 dvss 0.0469527
R13625 dvss.n2815 dvss 0.0469527
R13626 dvss.n2768 dvss 0.0469527
R13627 dvss.n2721 dvss 0.0469527
R13628 dvss.n2674 dvss 0.0469527
R13629 dvss.n2627 dvss 0.0469527
R13630 dvss.n2927 dvss 0.0469527
R13631 dvss.n2285 dvss 0.0469527
R13632 dvss.n4112 dvss 0.0469527
R13633 dvss.n4065 dvss 0.0469527
R13634 dvss dvss.n2834 0.0435743
R13635 dvss.n2823 dvss 0.0435743
R13636 dvss dvss.n2787 0.0435743
R13637 dvss.n2776 dvss 0.0435743
R13638 dvss dvss.n2740 0.0435743
R13639 dvss.n2729 dvss 0.0435743
R13640 dvss dvss.n2693 0.0435743
R13641 dvss.n2682 dvss 0.0435743
R13642 dvss dvss.n2646 0.0435743
R13643 dvss.n2635 dvss 0.0435743
R13644 dvss.n2905 dvss 0.0435743
R13645 dvss dvss.n2310 0.0435743
R13646 dvss.n2980 dvss 0.0435743
R13647 dvss.n2231 dvss 0.0435743
R13648 dvss.n4116 dvss 0.0435743
R13649 dvss dvss.n363 0.0435743
R13650 dvss dvss.n4084 0.0435743
R13651 dvss.n4073 dvss 0.0435743
R13652 dvss dvss.n2855 0.0410405
R13653 dvss.n2426 dvss 0.0410405
R13654 dvss.n2806 dvss 0.0410405
R13655 dvss.n2459 dvss 0.0410405
R13656 dvss.n2759 dvss 0.0410405
R13657 dvss.n2495 dvss 0.0410405
R13658 dvss.n2712 dvss 0.0410405
R13659 dvss.n2531 dvss 0.0410405
R13660 dvss.n2665 dvss 0.0410405
R13661 dvss.n2567 dvss 0.0410405
R13662 dvss.n2618 dvss 0.0410405
R13663 dvss.n2603 dvss 0.0410405
R13664 dvss dvss.n2941 0.0410405
R13665 dvss dvss.n2298 0.0410405
R13666 dvss.n2276 dvss 0.0410405
R13667 dvss.n2271 dvss 0.0410405
R13668 dvss.n4103 dvss 0.0410405
R13669 dvss.n281 dvss 0.0410405
R13670 dvss dvss.n2862 0.0385068
R13671 dvss.n4039 dvss.n4038 0.0362143
R13672 dvss dvss.n2859 0.0351284
R13673 dvss.n1059 dvss 0.0323548
R13674 dvss.n1060 dvss 0.0323548
R13675 dvss.n1065 dvss 0.0323548
R13676 dvss.n1066 dvss 0.0323548
R13677 dvss.n1067 dvss 0.0323548
R13678 dvss.n1068 dvss 0.0323548
R13679 dvss.n1078 dvss 0.0323548
R13680 dvss.n1079 dvss 0.0323548
R13681 dvss.n1090 dvss 0.0323548
R13682 dvss.n1091 dvss 0.0323548
R13683 dvss.n1103 dvss 0.0323548
R13684 dvss.n1105 dvss 0.0323548
R13685 dvss.n1109 dvss 0.0323548
R13686 dvss.n1110 dvss 0.0323548
R13687 dvss.n1133 dvss 0.0323548
R13688 dvss.n1119 dvss 0.0323548
R13689 dvss.n1146 dvss 0.0323548
R13690 dvss.n1147 dvss 0.0323548
R13691 dvss.n1162 dvss 0.0323548
R13692 dvss dvss.n1161 0.0323548
R13693 dvss.n1497 dvss 0.0323548
R13694 dvss.n1498 dvss 0.0323548
R13695 dvss.n1500 dvss 0.0323548
R13696 dvss dvss.n1499 0.0323548
R13697 dvss.n1509 dvss 0.0323548
R13698 dvss.n1512 dvss 0.0323548
R13699 dvss dvss.n1511 0.0323548
R13700 dvss.n1527 dvss 0.0323548
R13701 dvss dvss.n832 0.0323548
R13702 dvss.n1551 dvss 0.0323548
R13703 dvss.n1552 dvss 0.0323548
R13704 dvss.n1565 dvss 0.0323548
R13705 dvss.n1566 dvss 0.0323548
R13706 dvss.n1670 dvss 0.0323548
R13707 dvss dvss.n1669 0.0323548
R13708 dvss dvss.n1668 0.0323548
R13709 dvss.n1665 dvss 0.0323548
R13710 dvss dvss.n1663 0.0323548
R13711 dvss.n1660 dvss 0.0323548
R13712 dvss dvss.n1659 0.0323548
R13713 dvss.n1651 dvss 0.0323548
R13714 dvss.n1642 dvss 0.0323548
R13715 dvss.n1634 dvss 0.0323548
R13716 dvss dvss.n1633 0.0323548
R13717 dvss.n1624 dvss 0.0323548
R13718 dvss dvss.n1623 0.0323548
R13719 dvss.n1972 dvss 0.0323548
R13720 dvss.n1973 dvss 0.0323548
R13721 dvss.n1975 dvss 0.0323548
R13722 dvss dvss.n1974 0.0323548
R13723 dvss.n1984 dvss 0.0323548
R13724 dvss.n1987 dvss 0.0323548
R13725 dvss dvss.n1986 0.0323548
R13726 dvss.n2002 dvss 0.0323548
R13727 dvss dvss.n723 0.0323548
R13728 dvss.n2026 dvss 0.0323548
R13729 dvss.n2027 dvss 0.0323548
R13730 dvss.n2040 dvss 0.0323548
R13731 dvss.n2041 dvss 0.0323548
R13732 dvss.n3148 dvss 0.0323548
R13733 dvss dvss.n3147 0.0323548
R13734 dvss dvss.n3146 0.0323548
R13735 dvss.n3143 dvss 0.0323548
R13736 dvss dvss.n3141 0.0323548
R13737 dvss.n3138 dvss 0.0323548
R13738 dvss dvss.n3137 0.0323548
R13739 dvss.n3129 dvss 0.0323548
R13740 dvss.n3120 dvss 0.0323548
R13741 dvss.n3112 dvss 0.0323548
R13742 dvss dvss.n3111 0.0323548
R13743 dvss.n3102 dvss 0.0323548
R13744 dvss dvss.n3101 0.0323548
R13745 dvss dvss.n3100 0.0323548
R13746 dvss.n3097 dvss 0.0323548
R13747 dvss dvss.n3096 0.0323548
R13748 dvss dvss.n3095 0.0323548
R13749 dvss dvss.n3091 0.0323548
R13750 dvss dvss.n3090 0.0323548
R13751 dvss.n3087 dvss 0.0323548
R13752 dvss.n3079 dvss 0.0323548
R13753 dvss.n3070 dvss 0.0323548
R13754 dvss.n3062 dvss 0.0323548
R13755 dvss dvss.n3061 0.0323548
R13756 dvss.n3052 dvss 0.0323548
R13757 dvss dvss.n3051 0.0323548
R13758 dvss dvss.n3050 0.0323548
R13759 dvss.n3047 dvss 0.0323548
R13760 dvss dvss.n3046 0.0323548
R13761 dvss dvss.n3045 0.0323548
R13762 dvss dvss.n3041 0.0323548
R13763 dvss dvss.n3040 0.0323548
R13764 dvss.n3037 dvss 0.0323548
R13765 dvss.n3029 dvss 0.0323548
R13766 dvss.n3020 dvss 0.0323548
R13767 dvss.n3012 dvss 0.0323548
R13768 dvss dvss.n3011 0.0323548
R13769 dvss.n3002 dvss 0.0323548
R13770 dvss dvss.n3001 0.0323548
R13771 dvss.n3630 dvss 0.0323548
R13772 dvss.n3631 dvss 0.0323548
R13773 dvss.n3633 dvss 0.0323548
R13774 dvss dvss.n3632 0.0323548
R13775 dvss.n3642 dvss 0.0323548
R13776 dvss.n3645 dvss 0.0323548
R13777 dvss dvss.n3644 0.0323548
R13778 dvss.n3660 dvss 0.0323548
R13779 dvss dvss.n487 0.0323548
R13780 dvss.n3684 dvss 0.0323548
R13781 dvss.n3685 dvss 0.0323548
R13782 dvss.n3698 dvss 0.0323548
R13783 dvss.n3699 dvss 0.0323548
R13784 dvss.n3805 dvss 0.0323548
R13785 dvss dvss.n3804 0.0323548
R13786 dvss dvss.n3803 0.0323548
R13787 dvss.n3800 dvss 0.0323548
R13788 dvss dvss.n3798 0.0323548
R13789 dvss.n3795 dvss 0.0323548
R13790 dvss dvss.n3794 0.0323548
R13791 dvss.n3786 dvss 0.0323548
R13792 dvss.n3777 dvss 0.0323548
R13793 dvss.n3769 dvss 0.0323548
R13794 dvss dvss.n3768 0.0323548
R13795 dvss.n3759 dvss 0.0323548
R13796 dvss dvss.n3758 0.0323548
R13797 dvss dvss.n3757 0.0323548
R13798 dvss.n4050 dvss 0.0323548
R13799 dvss dvss.n4049 0.0323548
R13800 dvss dvss.n4048 0.0323548
R13801 dvss.n1142 dvss 0.0319516
R13802 dvss dvss.n828 0.0319516
R13803 dvss dvss.n1641 0.0319516
R13804 dvss dvss.n719 0.0319516
R13805 dvss dvss.n3119 0.0319516
R13806 dvss dvss.n3069 0.0319516
R13807 dvss dvss.n3019 0.0319516
R13808 dvss dvss.n483 0.0319516
R13809 dvss dvss.n3776 0.0319516
R13810 dvss.n4021 dvss.n4015 0.0310921
R13811 dvss.n4028 dvss.n4024 0.0310921
R13812 dvss dvss.n2830 0.0300608
R13813 dvss dvss.n2783 0.0300608
R13814 dvss dvss.n2736 0.0300608
R13815 dvss dvss.n2689 0.0300608
R13816 dvss dvss.n2642 0.0300608
R13817 dvss.n2909 dvss 0.0300608
R13818 dvss.n2223 dvss 0.0300608
R13819 dvss.n358 dvss 0.0300608
R13820 dvss dvss.n4080 0.0300608
R13821 dvss.n1074 dvss 0.0287258
R13822 dvss.n1238 dvss 0.0282388
R13823 dvss.n1264 dvss 0.0282388
R13824 dvss dvss.n1275 0.0282388
R13825 dvss dvss.n1302 0.0282388
R13826 dvss dvss.n1316 0.0282388
R13827 dvss.n1326 dvss 0.0282388
R13828 dvss.n1484 dvss 0.0282388
R13829 dvss dvss.n1483 0.0282388
R13830 dvss dvss.n1482 0.0282388
R13831 dvss dvss.n1478 0.0282388
R13832 dvss.n1410 dvss 0.0282388
R13833 dvss dvss.n1461 0.0282388
R13834 dvss dvss.n1450 0.0282388
R13835 dvss.n1437 dvss 0.0282388
R13836 dvss.n1679 dvss 0.0282388
R13837 dvss.n1704 dvss 0.0282388
R13838 dvss.n1701 dvss 0.0282388
R13839 dvss dvss.n1700 0.0282388
R13840 dvss.n1713 dvss 0.0282388
R13841 dvss.n1739 dvss 0.0282388
R13842 dvss dvss.n1750 0.0282388
R13843 dvss dvss.n1777 0.0282388
R13844 dvss dvss.n1791 0.0282388
R13845 dvss.n1801 dvss 0.0282388
R13846 dvss.n1959 dvss 0.0282388
R13847 dvss dvss.n1958 0.0282388
R13848 dvss dvss.n1957 0.0282388
R13849 dvss dvss.n1953 0.0282388
R13850 dvss.n1885 dvss 0.0282388
R13851 dvss dvss.n1936 0.0282388
R13852 dvss dvss.n1925 0.0282388
R13853 dvss.n1912 dvss 0.0282388
R13854 dvss.n3157 dvss 0.0282388
R13855 dvss.n3182 dvss 0.0282388
R13856 dvss.n3179 dvss 0.0282388
R13857 dvss dvss.n3178 0.0282388
R13858 dvss.n3191 dvss 0.0282388
R13859 dvss.n3217 dvss 0.0282388
R13860 dvss dvss.n3228 0.0282388
R13861 dvss dvss.n3255 0.0282388
R13862 dvss dvss.n3270 0.0282388
R13863 dvss.n3280 dvss 0.0282388
R13864 dvss dvss.n642 0.0282388
R13865 dvss.n3302 dvss 0.0282388
R13866 dvss.n3299 dvss 0.0282388
R13867 dvss.n3310 dvss 0.0282388
R13868 dvss.n3342 dvss 0.0282388
R13869 dvss.n3354 dvss 0.0282388
R13870 dvss.n3376 dvss 0.0282388
R13871 dvss dvss.n3387 0.0282388
R13872 dvss.n3397 dvss 0.0282388
R13873 dvss dvss.n3400 0.0282388
R13874 dvss.n3415 dvss 0.0282388
R13875 dvss dvss.n3414 0.0282388
R13876 dvss.n3423 dvss 0.0282388
R13877 dvss.n3449 dvss 0.0282388
R13878 dvss dvss.n3457 0.0282388
R13879 dvss dvss.n3487 0.0282388
R13880 dvss dvss.n3501 0.0282388
R13881 dvss.n3511 dvss 0.0282388
R13882 dvss.n3617 dvss 0.0282388
R13883 dvss dvss.n3616 0.0282388
R13884 dvss dvss.n3615 0.0282388
R13885 dvss dvss.n3611 0.0282388
R13886 dvss.n3550 dvss 0.0282388
R13887 dvss dvss.n3594 0.0282388
R13888 dvss dvss.n3888 0.0282388
R13889 dvss.n460 dvss 0.0282388
R13890 dvss.n461 dvss 0.0282388
R13891 dvss.n3873 dvss 0.0282388
R13892 dvss dvss.n3872 0.0282388
R13893 dvss dvss.n3871 0.0282388
R13894 dvss dvss.n3867 0.0282388
R13895 dvss.n3828 dvss 0.0282388
R13896 dvss dvss.n3850 0.0282388
R13897 dvss.n3946 dvss 0.0282388
R13898 dvss.n3963 dvss 0.0282388
R13899 dvss dvss.n3962 0.0282388
R13900 dvss.n3977 dvss 0.0282388
R13901 dvss.n3978 dvss 0.0282388
R13902 dvss.n3985 dvss 0.0282388
R13903 dvss.n961 dvss 0.0278876
R13904 dvss.n959 dvss 0.0278876
R13905 dvss.n970 dvss 0.0278876
R13906 dvss.n972 dvss 0.0278876
R13907 dvss.n974 dvss 0.0278876
R13908 dvss.n956 dvss 0.0278876
R13909 dvss.n989 dvss 0.0278876
R13910 dvss.n953 dvss 0.0278876
R13911 dvss.n1009 dvss 0.0278876
R13912 dvss.n1011 dvss 0.0278876
R13913 dvss.n939 dvss 0.0278876
R13914 dvss.n1289 dvss 0.0278876
R13915 dvss dvss.n1460 0.0278876
R13916 dvss.n1764 dvss 0.0278876
R13917 dvss dvss.n1935 0.0278876
R13918 dvss.n3242 dvss 0.0278876
R13919 dvss.n3358 dvss 0.0278876
R13920 dvss.n3474 dvss 0.0278876
R13921 dvss dvss.n3593 0.0278876
R13922 dvss dvss.n3849 0.0278876
R13923 dvss.n1244 dvss 0.0257809
R13924 dvss dvss.n1474 0.0257809
R13925 dvss.n1719 dvss 0.0257809
R13926 dvss dvss.n1949 0.0257809
R13927 dvss.n3197 dvss 0.0257809
R13928 dvss.n3319 dvss 0.0257809
R13929 dvss.n3438 dvss 0.0257809
R13930 dvss dvss.n3607 0.0257809
R13931 dvss dvss.n3863 0.0257809
R13932 dvss.n984 dvss 0.0247275
R13933 dvss.n2831 dvss 0.0233041
R13934 dvss.n2784 dvss 0.0233041
R13935 dvss.n2737 dvss 0.0233041
R13936 dvss.n2690 dvss 0.0233041
R13937 dvss.n2643 dvss 0.0233041
R13938 dvss.n2907 dvss 0.0233041
R13939 dvss dvss.n2982 0.0233041
R13940 dvss dvss.n4118 0.0233041
R13941 dvss.n4081 dvss 0.0233041
R13942 dvss dvss.n1112 0.0230806
R13943 dvss dvss.n1521 0.0230806
R13944 dvss dvss.n1654 0.0230806
R13945 dvss dvss.n1996 0.0230806
R13946 dvss dvss.n3132 0.0230806
R13947 dvss dvss.n3082 0.0230806
R13948 dvss dvss.n3032 0.0230806
R13949 dvss dvss.n3654 0.0230806
R13950 dvss dvss.n3789 0.0230806
R13951 dvss.n1088 dvss 0.0226774
R13952 dvss.n1159 dvss 0.0226774
R13953 dvss.n822 dvss 0.0226774
R13954 dvss dvss.n1628 0.0226774
R13955 dvss.n713 dvss 0.0226774
R13956 dvss dvss.n3106 0.0226774
R13957 dvss dvss.n3056 0.0226774
R13958 dvss dvss.n3006 0.0226774
R13959 dvss.n477 dvss 0.0226774
R13960 dvss dvss.n3763 0.0226774
R13961 dvss.n143 dvss 0.0226354
R13962 dvss dvss.n153 0.0226354
R13963 dvss.n246 dvss 0.0226354
R13964 dvss dvss.n256 0.0226354
R13965 dvss.n164 dvss 0.0226354
R13966 dvss.n155 dvss 0.0226354
R13967 dvss.n228 dvss 0.0226354
R13968 dvss dvss.n0 0.0226354
R13969 dvss.n4136 dvss 0.0226354
R13970 dvss.n1134 dvss 0.0222742
R13971 dvss.n1144 dvss 0.0222742
R13972 dvss dvss.n1526 0.0222742
R13973 dvss dvss.n1541 0.0222742
R13974 dvss dvss.n1650 0.0222742
R13975 dvss.n1638 dvss 0.0222742
R13976 dvss dvss.n2001 0.0222742
R13977 dvss dvss.n2016 0.0222742
R13978 dvss dvss.n3128 0.0222742
R13979 dvss.n3116 dvss 0.0222742
R13980 dvss dvss.n3078 0.0222742
R13981 dvss.n3066 dvss 0.0222742
R13982 dvss dvss.n3028 0.0222742
R13983 dvss.n3016 dvss 0.0222742
R13984 dvss dvss.n3659 0.0222742
R13985 dvss dvss.n3674 0.0222742
R13986 dvss dvss.n3785 0.0222742
R13987 dvss.n3773 dvss 0.0222742
R13988 dvss.n1154 dvss 0.0202581
R13989 dvss.n1557 dvss 0.0202581
R13990 dvss.n1591 dvss 0.0202581
R13991 dvss.n2032 dvss 0.0202581
R13992 dvss.n2066 dvss 0.0202581
R13993 dvss.n2097 dvss 0.0202581
R13994 dvss.n2128 dvss 0.0202581
R13995 dvss.n3690 dvss 0.0202581
R13996 dvss.n3740 dvss 0.0202581
R13997 dvss.n1257 dvss 0.0201629
R13998 dvss.n1409 dvss 0.0201629
R13999 dvss.n1732 dvss 0.0201629
R14000 dvss.n1884 dvss 0.0201629
R14001 dvss.n3210 dvss 0.0201629
R14002 dvss dvss.n3330 0.0201629
R14003 dvss.n3448 dvss 0.0201629
R14004 dvss.n3549 dvss 0.0201629
R14005 dvss.n3827 dvss 0.0201629
R14006 dvss.n1508 dvss 0.0198548
R14007 dvss dvss.n1664 0.0198548
R14008 dvss.n1983 dvss 0.0198548
R14009 dvss dvss.n3142 0.0198548
R14010 dvss.n3092 dvss 0.0198548
R14011 dvss.n3042 dvss 0.0198548
R14012 dvss.n3641 dvss 0.0198548
R14013 dvss dvss.n3799 0.0198548
R14014 dvss dvss.n860 0.0198118
R14015 dvss.n1682 dvss 0.0198118
R14016 dvss dvss.n751 0.0198118
R14017 dvss.n3160 dvss 0.0198118
R14018 dvss dvss.n641 0.0198118
R14019 dvss dvss.n579 0.0198118
R14020 dvss dvss.n516 0.0198118
R14021 dvss.n3877 dvss 0.0198118
R14022 dvss dvss.n322 0.0198118
R14023 dvss.n1265 dvss 0.0194607
R14024 dvss.n1466 dvss 0.0194607
R14025 dvss.n1740 dvss 0.0194607
R14026 dvss.n1941 dvss 0.0194607
R14027 dvss.n3218 dvss 0.0194607
R14028 dvss dvss.n3341 0.0194607
R14029 dvss.n3450 dvss 0.0194607
R14030 dvss.n3599 dvss 0.0194607
R14031 dvss.n3855 dvss 0.0194607
R14032 dvss.n1104 dvss 0.0194516
R14033 dvss.n1076 dvss 0.0190484
R14034 dvss.n1099 dvss 0.0186452
R14035 dvss dvss.n881 0.0184073
R14036 dvss.n1359 dvss 0.0184073
R14037 dvss dvss.n772 0.0184073
R14038 dvss.n1834 dvss 0.0184073
R14039 dvss dvss.n663 0.0184073
R14040 dvss dvss.n603 0.0184073
R14041 dvss dvss.n537 0.0184073
R14042 dvss.n3587 dvss 0.0184073
R14043 dvss.n3843 dvss 0.0184073
R14044 dvss.n2860 dvss 0.0182365
R14045 dvss dvss.n901 0.0173539
R14046 dvss.n1479 dvss 0.0173539
R14047 dvss.n1339 dvss 0.0173539
R14048 dvss dvss.n1699 0.0173539
R14049 dvss dvss.n792 0.0173539
R14050 dvss.n1954 dvss 0.0173539
R14051 dvss.n1814 dvss 0.0173539
R14052 dvss dvss.n3177 0.0173539
R14053 dvss dvss.n683 0.0173539
R14054 dvss dvss.n3298 0.0173539
R14055 dvss.n3316 dvss 0.0173539
R14056 dvss dvss.n3413 0.0173539
R14057 dvss.n3429 dvss 0.0173539
R14058 dvss.n3612 dvss 0.0173539
R14059 dvss.n3524 dvss 0.0173539
R14060 dvss.n3868 dvss 0.0173539
R14061 dvss.n403 dvss 0.0173539
R14062 dvss.n1102 dvss 0.0170323
R14063 dvss.n948 dvss 0.0170028
R14064 dvss dvss.n997 0.0166517
R14065 dvss.n986 dvss 0.0163006
R14066 dvss.n1321 dvss 0.0163006
R14067 dvss dvss.n865 0.0163006
R14068 dvss.n1443 dvss 0.0163006
R14069 dvss dvss.n1445 0.0163006
R14070 dvss.n1796 dvss 0.0163006
R14071 dvss dvss.n756 0.0163006
R14072 dvss.n1918 dvss 0.0163006
R14073 dvss dvss.n1920 0.0163006
R14074 dvss.n3275 dvss 0.0163006
R14075 dvss dvss.n647 0.0163006
R14076 dvss.n3392 dvss 0.0163006
R14077 dvss dvss.n584 0.0163006
R14078 dvss.n3506 dvss 0.0163006
R14079 dvss dvss.n521 0.0163006
R14080 dvss.n3881 dvss 0.0163006
R14081 dvss dvss.n3883 0.0163006
R14082 dvss.n3957 dvss 0.0163006
R14083 dvss dvss.n336 0.0163006
R14084 dvss.n1026 dvss 0.0159494
R14085 dvss.n2886 dvss 0.0148581
R14086 dvss.n2885 dvss 0.0148581
R14087 dvss.n2882 dvss 0.0148581
R14088 dvss.n2881 dvss 0.0148581
R14089 dvss.n2880 dvss 0.0148581
R14090 dvss.n2877 dvss 0.0148581
R14091 dvss.n2876 dvss 0.0148581
R14092 dvss.n2875 dvss 0.0148581
R14093 dvss.n2872 dvss 0.0148581
R14094 dvss.n2871 dvss 0.0148581
R14095 dvss.n2870 dvss 0.0148581
R14096 dvss.n2864 dvss 0.0148581
R14097 dvss.n2863 dvss 0.0148581
R14098 dvss.n2862 dvss 0.0148581
R14099 dvss.n2415 dvss 0.0148581
R14100 dvss.n2415 dvss 0.0148581
R14101 dvss.n2860 dvss 0.0148581
R14102 dvss.n2859 dvss 0.0148581
R14103 dvss.n2856 dvss 0.0148581
R14104 dvss.n2855 dvss 0.0148581
R14105 dvss.n2852 dvss 0.0148581
R14106 dvss.n2851 dvss 0.0148581
R14107 dvss.n2848 dvss 0.0148581
R14108 dvss.n2845 dvss 0.0148581
R14109 dvss.n2844 dvss 0.0148581
R14110 dvss.n2843 dvss 0.0148581
R14111 dvss.n2840 dvss 0.0148581
R14112 dvss.n2839 dvss 0.0148581
R14113 dvss.n2838 dvss 0.0148581
R14114 dvss.n2835 dvss 0.0148581
R14115 dvss.n2834 dvss 0.0148581
R14116 dvss dvss.n2439 0.0148581
R14117 dvss.n2831 dvss 0.0148581
R14118 dvss.n2830 dvss 0.0148581
R14119 dvss.n2827 dvss 0.0148581
R14120 dvss.n2823 dvss 0.0148581
R14121 dvss.n2822 dvss 0.0148581
R14122 dvss.n2819 dvss 0.0148581
R14123 dvss.n2818 dvss 0.0148581
R14124 dvss.n2817 dvss 0.0148581
R14125 dvss.n2811 dvss 0.0148581
R14126 dvss.n2810 dvss 0.0148581
R14127 dvss.n2809 dvss 0.0148581
R14128 dvss.n2806 dvss 0.0148581
R14129 dvss.n2805 dvss 0.0148581
R14130 dvss.n2804 dvss 0.0148581
R14131 dvss.n2801 dvss 0.0148581
R14132 dvss.n2798 dvss 0.0148581
R14133 dvss.n2797 dvss 0.0148581
R14134 dvss.n2796 dvss 0.0148581
R14135 dvss.n2793 dvss 0.0148581
R14136 dvss.n2792 dvss 0.0148581
R14137 dvss.n2791 dvss 0.0148581
R14138 dvss.n2788 dvss 0.0148581
R14139 dvss.n2787 dvss 0.0148581
R14140 dvss dvss.n2475 0.0148581
R14141 dvss.n2784 dvss 0.0148581
R14142 dvss.n2783 dvss 0.0148581
R14143 dvss.n2780 dvss 0.0148581
R14144 dvss.n2776 dvss 0.0148581
R14145 dvss.n2775 dvss 0.0148581
R14146 dvss.n2772 dvss 0.0148581
R14147 dvss.n2771 dvss 0.0148581
R14148 dvss.n2770 dvss 0.0148581
R14149 dvss.n2764 dvss 0.0148581
R14150 dvss.n2763 dvss 0.0148581
R14151 dvss.n2762 dvss 0.0148581
R14152 dvss.n2759 dvss 0.0148581
R14153 dvss.n2758 dvss 0.0148581
R14154 dvss.n2757 dvss 0.0148581
R14155 dvss.n2754 dvss 0.0148581
R14156 dvss.n2751 dvss 0.0148581
R14157 dvss.n2750 dvss 0.0148581
R14158 dvss.n2749 dvss 0.0148581
R14159 dvss.n2746 dvss 0.0148581
R14160 dvss.n2745 dvss 0.0148581
R14161 dvss.n2744 dvss 0.0148581
R14162 dvss.n2741 dvss 0.0148581
R14163 dvss.n2740 dvss 0.0148581
R14164 dvss dvss.n2511 0.0148581
R14165 dvss.n2737 dvss 0.0148581
R14166 dvss.n2736 dvss 0.0148581
R14167 dvss.n2733 dvss 0.0148581
R14168 dvss.n2729 dvss 0.0148581
R14169 dvss.n2728 dvss 0.0148581
R14170 dvss.n2725 dvss 0.0148581
R14171 dvss.n2724 dvss 0.0148581
R14172 dvss.n2723 dvss 0.0148581
R14173 dvss.n2717 dvss 0.0148581
R14174 dvss.n2716 dvss 0.0148581
R14175 dvss.n2715 dvss 0.0148581
R14176 dvss.n2712 dvss 0.0148581
R14177 dvss.n2711 dvss 0.0148581
R14178 dvss.n2710 dvss 0.0148581
R14179 dvss.n2707 dvss 0.0148581
R14180 dvss.n2704 dvss 0.0148581
R14181 dvss.n2703 dvss 0.0148581
R14182 dvss.n2702 dvss 0.0148581
R14183 dvss.n2699 dvss 0.0148581
R14184 dvss.n2698 dvss 0.0148581
R14185 dvss.n2697 dvss 0.0148581
R14186 dvss.n2694 dvss 0.0148581
R14187 dvss.n2693 dvss 0.0148581
R14188 dvss dvss.n2547 0.0148581
R14189 dvss.n2690 dvss 0.0148581
R14190 dvss.n2689 dvss 0.0148581
R14191 dvss.n2686 dvss 0.0148581
R14192 dvss.n2682 dvss 0.0148581
R14193 dvss.n2681 dvss 0.0148581
R14194 dvss.n2678 dvss 0.0148581
R14195 dvss.n2677 dvss 0.0148581
R14196 dvss.n2676 dvss 0.0148581
R14197 dvss.n2670 dvss 0.0148581
R14198 dvss.n2669 dvss 0.0148581
R14199 dvss.n2668 dvss 0.0148581
R14200 dvss.n2665 dvss 0.0148581
R14201 dvss.n2664 dvss 0.0148581
R14202 dvss.n2663 dvss 0.0148581
R14203 dvss.n2660 dvss 0.0148581
R14204 dvss.n2657 dvss 0.0148581
R14205 dvss.n2656 dvss 0.0148581
R14206 dvss.n2655 dvss 0.0148581
R14207 dvss.n2652 dvss 0.0148581
R14208 dvss.n2651 dvss 0.0148581
R14209 dvss.n2650 dvss 0.0148581
R14210 dvss.n2647 dvss 0.0148581
R14211 dvss.n2646 dvss 0.0148581
R14212 dvss dvss.n2583 0.0148581
R14213 dvss.n2643 dvss 0.0148581
R14214 dvss.n2642 dvss 0.0148581
R14215 dvss.n2639 dvss 0.0148581
R14216 dvss.n2635 dvss 0.0148581
R14217 dvss.n2634 dvss 0.0148581
R14218 dvss.n2631 dvss 0.0148581
R14219 dvss.n2630 dvss 0.0148581
R14220 dvss.n2629 dvss 0.0148581
R14221 dvss.n2623 dvss 0.0148581
R14222 dvss.n2622 dvss 0.0148581
R14223 dvss.n2621 dvss 0.0148581
R14224 dvss.n2618 dvss 0.0148581
R14225 dvss.n2617 dvss 0.0148581
R14226 dvss.n2616 dvss 0.0148581
R14227 dvss.n2613 dvss 0.0148581
R14228 dvss.n2610 dvss 0.0148581
R14229 dvss.n2609 dvss 0.0148581
R14230 dvss dvss.n2893 0.0148581
R14231 dvss dvss.n2894 0.0148581
R14232 dvss.n2896 dvss 0.0148581
R14233 dvss.n2895 dvss 0.0148581
R14234 dvss dvss.n2904 0.0148581
R14235 dvss dvss.n2905 0.0148581
R14236 dvss dvss.n2906 0.0148581
R14237 dvss dvss.n2907 0.0148581
R14238 dvss.n2909 dvss 0.0148581
R14239 dvss.n2908 dvss 0.0148581
R14240 dvss dvss.n2310 0.0148581
R14241 dvss.n2919 dvss 0.0148581
R14242 dvss.n2918 dvss 0.0148581
R14243 dvss.n2930 dvss 0.0148581
R14244 dvss.n2929 dvss 0.0148581
R14245 dvss dvss.n2939 0.0148581
R14246 dvss dvss.n2940 0.0148581
R14247 dvss.n2942 dvss 0.0148581
R14248 dvss.n2941 dvss 0.0148581
R14249 dvss dvss.n2951 0.0148581
R14250 dvss.n2952 dvss 0.0148581
R14251 dvss.n2958 dvss 0.0148581
R14252 dvss.n2957 dvss 0.0148581
R14253 dvss dvss.n2966 0.0148581
R14254 dvss dvss.n2967 0.0148581
R14255 dvss.n2969 dvss 0.0148581
R14256 dvss.n2968 dvss 0.0148581
R14257 dvss dvss.n2978 0.0148581
R14258 dvss dvss.n2979 0.0148581
R14259 dvss.n2980 dvss 0.0148581
R14260 dvss.n2983 dvss 0.0148581
R14261 dvss.n2982 dvss 0.0148581
R14262 dvss dvss.n2223 0.0148581
R14263 dvss dvss.n2228 0.0148581
R14264 dvss dvss.n2231 0.0148581
R14265 dvss.n2234 dvss 0.0148581
R14266 dvss.n2233 dvss 0.0148581
R14267 dvss.n2232 dvss 0.0148581
R14268 dvss dvss.n2216 0.0148581
R14269 dvss.n2281 dvss 0.0148581
R14270 dvss.n2280 dvss 0.0148581
R14271 dvss.n2279 dvss 0.0148581
R14272 dvss.n2276 dvss 0.0148581
R14273 dvss.n2275 dvss 0.0148581
R14274 dvss.n2274 dvss 0.0148581
R14275 dvss.n4132 dvss 0.0148581
R14276 dvss.n4129 dvss 0.0148581
R14277 dvss.n4128 dvss 0.0148581
R14278 dvss.n4127 dvss 0.0148581
R14279 dvss.n4124 dvss 0.0148581
R14280 dvss.n4123 dvss 0.0148581
R14281 dvss.n4122 dvss 0.0148581
R14282 dvss.n4116 dvss 0.0148581
R14283 dvss.n4119 dvss 0.0148581
R14284 dvss.n4118 dvss 0.0148581
R14285 dvss dvss.n358 0.0148581
R14286 dvss.n366 dvss 0.0148581
R14287 dvss.n363 dvss 0.0148581
R14288 dvss.n362 dvss 0.0148581
R14289 dvss.n360 dvss 0.0148581
R14290 dvss.n359 dvss 0.0148581
R14291 dvss dvss.n271 0.0148581
R14292 dvss.n4108 dvss 0.0148581
R14293 dvss.n4107 dvss 0.0148581
R14294 dvss.n4106 dvss 0.0148581
R14295 dvss.n4103 dvss 0.0148581
R14296 dvss.n4102 dvss 0.0148581
R14297 dvss.n4101 dvss 0.0148581
R14298 dvss.n4098 dvss 0.0148581
R14299 dvss.n4095 dvss 0.0148581
R14300 dvss.n4094 dvss 0.0148581
R14301 dvss.n4093 dvss 0.0148581
R14302 dvss.n4090 dvss 0.0148581
R14303 dvss.n4089 dvss 0.0148581
R14304 dvss.n4088 dvss 0.0148581
R14305 dvss.n4085 dvss 0.0148581
R14306 dvss.n4084 dvss 0.0148581
R14307 dvss dvss.n293 0.0148581
R14308 dvss.n4081 dvss 0.0148581
R14309 dvss.n4080 dvss 0.0148581
R14310 dvss.n4077 dvss 0.0148581
R14311 dvss.n4073 dvss 0.0148581
R14312 dvss.n4072 dvss 0.0148581
R14313 dvss.n4069 dvss 0.0148581
R14314 dvss.n4068 dvss 0.0148581
R14315 dvss.n4067 dvss 0.0148581
R14316 dvss.n4061 dvss 0.0148581
R14317 dvss.n4060 dvss 0.0148581
R14318 dvss.n4059 dvss 0.0148581
R14319 dvss dvss.n1018 0.0145449
R14320 dvss.n2867 dvss 0.0140135
R14321 dvss dvss.n1111 0.0134032
R14322 dvss dvss.n1118 0.0134032
R14323 dvss.n1520 dvss 0.0134032
R14324 dvss dvss.n1536 0.0134032
R14325 dvss.n1574 dvss 0.0134032
R14326 dvss dvss.n1645 0.0134032
R14327 dvss.n1995 dvss 0.0134032
R14328 dvss dvss.n2011 0.0134032
R14329 dvss.n2049 dvss 0.0134032
R14330 dvss dvss.n3123 0.0134032
R14331 dvss.n2081 dvss 0.0134032
R14332 dvss dvss.n3073 0.0134032
R14333 dvss.n2112 dvss 0.0134032
R14334 dvss dvss.n3023 0.0134032
R14335 dvss.n3653 dvss 0.0134032
R14336 dvss dvss.n3669 0.0134032
R14337 dvss.n3707 dvss 0.0134032
R14338 dvss dvss.n3780 0.0134032
R14339 dvss.n1303 dvss 0.0127893
R14340 dvss.n1451 dvss 0.0127893
R14341 dvss.n1778 dvss 0.0127893
R14342 dvss.n1926 dvss 0.0127893
R14343 dvss.n3256 dvss 0.0127893
R14344 dvss.n3369 dvss 0.0127893
R14345 dvss.n3488 dvss 0.0127893
R14346 dvss.n3889 dvss 0.0127893
R14347 dvss.n3937 dvss 0.0127893
R14348 dvss.n1127 dvss 0.0125968
R14349 dvss.n1138 dvss 0.0125968
R14350 dvss dvss.n1510 0.0125968
R14351 dvss.n1537 dvss 0.0125968
R14352 dvss dvss.n1658 0.0125968
R14353 dvss.n1646 dvss 0.0125968
R14354 dvss dvss.n1985 0.0125968
R14355 dvss.n2012 dvss 0.0125968
R14356 dvss dvss.n3136 0.0125968
R14357 dvss.n3124 dvss 0.0125968
R14358 dvss dvss.n3086 0.0125968
R14359 dvss.n3074 dvss 0.0125968
R14360 dvss dvss.n3036 0.0125968
R14361 dvss.n3024 dvss 0.0125968
R14362 dvss dvss.n3643 0.0125968
R14363 dvss.n3670 dvss 0.0125968
R14364 dvss dvss.n3793 0.0125968
R14365 dvss.n3781 dvss 0.0125968
R14366 dvss dvss.n2851 0.0123243
R14367 dvss dvss.n2804 0.0123243
R14368 dvss dvss.n2757 0.0123243
R14369 dvss dvss.n2710 0.0123243
R14370 dvss dvss.n2663 0.0123243
R14371 dvss dvss.n2616 0.0123243
R14372 dvss.n2952 dvss 0.0123243
R14373 dvss dvss.n2274 0.0123243
R14374 dvss dvss.n4101 0.0123243
R14375 dvss dvss.n1251 0.011736
R14376 dvss.n1276 dvss 0.011736
R14377 dvss.n1471 dvss 0.011736
R14378 dvss.n1462 dvss 0.011736
R14379 dvss dvss.n1726 0.011736
R14380 dvss.n1751 dvss 0.011736
R14381 dvss.n1946 dvss 0.011736
R14382 dvss.n1937 dvss 0.011736
R14383 dvss dvss.n3204 0.011736
R14384 dvss.n3229 dvss 0.011736
R14385 dvss dvss.n624 0.011736
R14386 dvss dvss.n3336 0.011736
R14387 dvss.n3433 dvss 0.011736
R14388 dvss.n3458 dvss 0.011736
R14389 dvss.n3604 dvss 0.011736
R14390 dvss.n3595 dvss 0.011736
R14391 dvss.n3860 dvss 0.011736
R14392 dvss.n3851 dvss 0.011736
R14393 dvss dvss.n2445 0.0114797
R14394 dvss.n2814 dvss 0.0114797
R14395 dvss dvss.n2481 0.0114797
R14396 dvss.n2767 dvss 0.0114797
R14397 dvss dvss.n2517 0.0114797
R14398 dvss.n2720 dvss 0.0114797
R14399 dvss dvss.n2553 0.0114797
R14400 dvss.n2673 dvss 0.0114797
R14401 dvss dvss.n2589 0.0114797
R14402 dvss.n2626 dvss 0.0114797
R14403 dvss.n2922 dvss 0.0114797
R14404 dvss.n2926 dvss 0.0114797
R14405 dvss dvss.n2230 0.0114797
R14406 dvss.n2284 dvss 0.0114797
R14407 dvss.n364 dvss 0.0114797
R14408 dvss.n4111 dvss 0.0114797
R14409 dvss dvss.n297 0.0114797
R14410 dvss.n4064 dvss 0.0114797
R14411 dvss.n1252 dvss 0.0110337
R14412 dvss dvss.n1271 0.0110337
R14413 dvss.n1346 dvss 0.0110337
R14414 dvss.n1456 dvss 0.0110337
R14415 dvss.n1727 dvss 0.0110337
R14416 dvss dvss.n1746 0.0110337
R14417 dvss.n1821 dvss 0.0110337
R14418 dvss.n1931 dvss 0.0110337
R14419 dvss.n3205 dvss 0.0110337
R14420 dvss dvss.n3224 0.0110337
R14421 dvss dvss.n625 0.0110337
R14422 dvss.n3337 dvss 0.0110337
R14423 dvss dvss.n3437 0.0110337
R14424 dvss.n3456 dvss 0.0110337
R14425 dvss.n3531 dvss 0.0110337
R14426 dvss.n3589 dvss 0.0110337
R14427 dvss.n410 dvss 0.0110337
R14428 dvss.n3845 dvss 0.0110337
R14429 dvss dvss.n1292 0.00998034
R14430 dvss.n1367 dvss 0.00998034
R14431 dvss dvss.n1767 0.00998034
R14432 dvss.n1842 dvss 0.00998034
R14433 dvss dvss.n3245 0.00998034
R14434 dvss dvss.n3361 0.00998034
R14435 dvss dvss.n3477 0.00998034
R14436 dvss.n384 dvss 0.00998034
R14437 dvss.n3936 dvss 0.00998034
R14438 dvss.n2439 dvss 0.00979054
R14439 dvss dvss.n2822 0.00979054
R14440 dvss.n2475 dvss 0.00979054
R14441 dvss dvss.n2775 0.00979054
R14442 dvss.n2511 dvss 0.00979054
R14443 dvss dvss.n2728 0.00979054
R14444 dvss.n2547 dvss 0.00979054
R14445 dvss dvss.n2681 0.00979054
R14446 dvss.n2583 dvss 0.00979054
R14447 dvss dvss.n2634 0.00979054
R14448 dvss.n2906 dvss 0.00979054
R14449 dvss.n2919 dvss 0.00979054
R14450 dvss.n2983 dvss 0.00979054
R14451 dvss.n2234 dvss 0.00979054
R14452 dvss.n4119 dvss 0.00979054
R14453 dvss dvss.n362 0.00979054
R14454 dvss.n293 dvss 0.00979054
R14455 dvss dvss.n4072 0.00979054
R14456 dvss.n1101 dvss 0.00896774
R14457 dvss.n2849 dvss 0.00894595
R14458 dvss.n2802 dvss 0.00894595
R14459 dvss.n2755 dvss 0.00894595
R14460 dvss.n2708 dvss 0.00894595
R14461 dvss.n2661 dvss 0.00894595
R14462 dvss.n2614 dvss 0.00894595
R14463 dvss dvss.n2956 0.00894595
R14464 dvss.n2272 dvss 0.00894595
R14465 dvss.n4099 dvss 0.00894595
R14466 dvss.n4133 dvss 0.00810135
R14467 dvss dvss.n1028 0.00752247
R14468 dvss dvss.n1059 0.00735484
R14469 dvss dvss.n1060 0.00735484
R14470 dvss dvss.n1065 0.00735484
R14471 dvss dvss.n1066 0.00735484
R14472 dvss dvss.n1067 0.00735484
R14473 dvss dvss.n1068 0.00735484
R14474 dvss dvss.n1076 0.00735484
R14475 dvss dvss.n1077 0.00735484
R14476 dvss dvss.n1078 0.00735484
R14477 dvss dvss.n1090 0.00735484
R14478 dvss dvss.n1091 0.00735484
R14479 dvss.n1099 dvss 0.00735484
R14480 dvss dvss.n1092 0.00735484
R14481 dvss dvss.n1092 0.00735484
R14482 dvss dvss.n1101 0.00735484
R14483 dvss dvss.n1102 0.00735484
R14484 dvss dvss.n1103 0.00735484
R14485 dvss dvss.n1104 0.00735484
R14486 dvss dvss.n1105 0.00735484
R14487 dvss dvss.n1109 0.00735484
R14488 dvss dvss.n1110 0.00735484
R14489 dvss.n1127 dvss 0.00735484
R14490 dvss dvss.n1111 0.00735484
R14491 dvss.n1130 dvss 0.00735484
R14492 dvss dvss.n1112 0.00735484
R14493 dvss dvss.n1133 0.00735484
R14494 dvss.n1134 dvss 0.00735484
R14495 dvss dvss.n1117 0.00735484
R14496 dvss.n1138 dvss 0.00735484
R14497 dvss dvss.n1118 0.00735484
R14498 dvss dvss.n1119 0.00735484
R14499 dvss dvss.n1144 0.00735484
R14500 dvss dvss.n1145 0.00735484
R14501 dvss dvss.n1146 0.00735484
R14502 dvss dvss.n1147 0.00735484
R14503 dvss dvss.n1152 0.00735484
R14504 dvss dvss.n1159 0.00735484
R14505 dvss dvss.n1160 0.00735484
R14506 dvss.n1162 dvss 0.00735484
R14507 dvss.n1161 dvss 0.00735484
R14508 dvss dvss.n1497 0.00735484
R14509 dvss dvss.n1498 0.00735484
R14510 dvss.n1500 dvss 0.00735484
R14511 dvss.n1499 dvss 0.00735484
R14512 dvss dvss.n1508 0.00735484
R14513 dvss dvss.n1509 0.00735484
R14514 dvss.n1512 dvss 0.00735484
R14515 dvss.n1511 dvss 0.00735484
R14516 dvss.n1510 dvss 0.00735484
R14517 dvss dvss.n1520 0.00735484
R14518 dvss.n1522 dvss 0.00735484
R14519 dvss.n1521 dvss 0.00735484
R14520 dvss.n1527 dvss 0.00735484
R14521 dvss.n1526 dvss 0.00735484
R14522 dvss.n838 dvss 0.00735484
R14523 dvss.n1537 dvss 0.00735484
R14524 dvss.n1536 dvss 0.00735484
R14525 dvss.n832 dvss 0.00735484
R14526 dvss.n1541 dvss 0.00735484
R14527 dvss.n829 dvss 0.00735484
R14528 dvss dvss.n1551 0.00735484
R14529 dvss dvss.n1552 0.00735484
R14530 dvss.n1553 dvss 0.00735484
R14531 dvss.n822 dvss 0.00735484
R14532 dvss.n821 dvss 0.00735484
R14533 dvss dvss.n1565 0.00735484
R14534 dvss dvss.n1566 0.00735484
R14535 dvss.n1670 dvss 0.00735484
R14536 dvss.n1669 dvss 0.00735484
R14537 dvss.n1668 dvss 0.00735484
R14538 dvss.n1665 dvss 0.00735484
R14539 dvss.n1664 dvss 0.00735484
R14540 dvss.n1663 dvss 0.00735484
R14541 dvss.n1660 dvss 0.00735484
R14542 dvss.n1659 dvss 0.00735484
R14543 dvss.n1658 dvss 0.00735484
R14544 dvss.n1574 dvss 0.00735484
R14545 dvss.n1655 dvss 0.00735484
R14546 dvss.n1654 dvss 0.00735484
R14547 dvss.n1651 dvss 0.00735484
R14548 dvss.n1650 dvss 0.00735484
R14549 dvss dvss.n1581 0.00735484
R14550 dvss.n1646 dvss 0.00735484
R14551 dvss.n1645 dvss 0.00735484
R14552 dvss.n1642 dvss 0.00735484
R14553 dvss.n1638 dvss 0.00735484
R14554 dvss.n1637 dvss 0.00735484
R14555 dvss.n1634 dvss 0.00735484
R14556 dvss.n1633 dvss 0.00735484
R14557 dvss.n1632 dvss 0.00735484
R14558 dvss.n1628 dvss 0.00735484
R14559 dvss.n1627 dvss 0.00735484
R14560 dvss.n1624 dvss 0.00735484
R14561 dvss.n1623 dvss 0.00735484
R14562 dvss dvss.n1972 0.00735484
R14563 dvss dvss.n1973 0.00735484
R14564 dvss.n1975 dvss 0.00735484
R14565 dvss.n1974 dvss 0.00735484
R14566 dvss dvss.n1983 0.00735484
R14567 dvss dvss.n1984 0.00735484
R14568 dvss.n1987 dvss 0.00735484
R14569 dvss.n1986 dvss 0.00735484
R14570 dvss.n1985 dvss 0.00735484
R14571 dvss dvss.n1995 0.00735484
R14572 dvss.n1997 dvss 0.00735484
R14573 dvss.n1996 dvss 0.00735484
R14574 dvss.n2002 dvss 0.00735484
R14575 dvss.n2001 dvss 0.00735484
R14576 dvss.n729 dvss 0.00735484
R14577 dvss.n2012 dvss 0.00735484
R14578 dvss.n2011 dvss 0.00735484
R14579 dvss.n723 dvss 0.00735484
R14580 dvss.n2016 dvss 0.00735484
R14581 dvss.n720 dvss 0.00735484
R14582 dvss dvss.n2026 0.00735484
R14583 dvss dvss.n2027 0.00735484
R14584 dvss.n2028 dvss 0.00735484
R14585 dvss.n713 dvss 0.00735484
R14586 dvss.n712 dvss 0.00735484
R14587 dvss dvss.n2040 0.00735484
R14588 dvss dvss.n2041 0.00735484
R14589 dvss.n3148 dvss 0.00735484
R14590 dvss.n3147 dvss 0.00735484
R14591 dvss.n3146 dvss 0.00735484
R14592 dvss.n3143 dvss 0.00735484
R14593 dvss.n3142 dvss 0.00735484
R14594 dvss.n3141 dvss 0.00735484
R14595 dvss.n3138 dvss 0.00735484
R14596 dvss.n3137 dvss 0.00735484
R14597 dvss.n3136 dvss 0.00735484
R14598 dvss.n2049 dvss 0.00735484
R14599 dvss.n3133 dvss 0.00735484
R14600 dvss.n3132 dvss 0.00735484
R14601 dvss.n3129 dvss 0.00735484
R14602 dvss.n3128 dvss 0.00735484
R14603 dvss dvss.n2056 0.00735484
R14604 dvss.n3124 dvss 0.00735484
R14605 dvss.n3123 dvss 0.00735484
R14606 dvss.n3120 dvss 0.00735484
R14607 dvss.n3116 dvss 0.00735484
R14608 dvss.n3115 dvss 0.00735484
R14609 dvss.n3112 dvss 0.00735484
R14610 dvss.n3111 dvss 0.00735484
R14611 dvss.n3110 dvss 0.00735484
R14612 dvss.n3106 dvss 0.00735484
R14613 dvss.n3105 dvss 0.00735484
R14614 dvss.n3102 dvss 0.00735484
R14615 dvss.n3101 dvss 0.00735484
R14616 dvss.n3100 dvss 0.00735484
R14617 dvss.n3097 dvss 0.00735484
R14618 dvss.n3096 dvss 0.00735484
R14619 dvss.n3095 dvss 0.00735484
R14620 dvss.n3092 dvss 0.00735484
R14621 dvss.n3091 dvss 0.00735484
R14622 dvss.n3090 dvss 0.00735484
R14623 dvss.n3087 dvss 0.00735484
R14624 dvss.n3086 dvss 0.00735484
R14625 dvss dvss.n2081 0.00735484
R14626 dvss.n3083 dvss 0.00735484
R14627 dvss.n3082 dvss 0.00735484
R14628 dvss.n3079 dvss 0.00735484
R14629 dvss.n3078 dvss 0.00735484
R14630 dvss dvss.n2087 0.00735484
R14631 dvss.n3074 dvss 0.00735484
R14632 dvss.n3073 dvss 0.00735484
R14633 dvss.n3070 dvss 0.00735484
R14634 dvss.n3066 dvss 0.00735484
R14635 dvss.n3065 dvss 0.00735484
R14636 dvss.n3062 dvss 0.00735484
R14637 dvss.n3061 dvss 0.00735484
R14638 dvss.n3060 dvss 0.00735484
R14639 dvss.n3056 dvss 0.00735484
R14640 dvss.n3055 dvss 0.00735484
R14641 dvss.n3052 dvss 0.00735484
R14642 dvss.n3051 dvss 0.00735484
R14643 dvss.n3050 dvss 0.00735484
R14644 dvss.n3047 dvss 0.00735484
R14645 dvss.n3046 dvss 0.00735484
R14646 dvss.n3045 dvss 0.00735484
R14647 dvss.n3042 dvss 0.00735484
R14648 dvss.n3041 dvss 0.00735484
R14649 dvss.n3040 dvss 0.00735484
R14650 dvss.n3037 dvss 0.00735484
R14651 dvss.n3036 dvss 0.00735484
R14652 dvss dvss.n2112 0.00735484
R14653 dvss.n3033 dvss 0.00735484
R14654 dvss.n3032 dvss 0.00735484
R14655 dvss.n3029 dvss 0.00735484
R14656 dvss.n3028 dvss 0.00735484
R14657 dvss dvss.n2118 0.00735484
R14658 dvss.n3024 dvss 0.00735484
R14659 dvss.n3023 dvss 0.00735484
R14660 dvss.n3020 dvss 0.00735484
R14661 dvss.n3016 dvss 0.00735484
R14662 dvss.n3015 dvss 0.00735484
R14663 dvss.n3012 dvss 0.00735484
R14664 dvss.n3011 dvss 0.00735484
R14665 dvss.n3010 dvss 0.00735484
R14666 dvss.n3006 dvss 0.00735484
R14667 dvss.n3005 dvss 0.00735484
R14668 dvss.n3002 dvss 0.00735484
R14669 dvss.n3001 dvss 0.00735484
R14670 dvss dvss.n3630 0.00735484
R14671 dvss dvss.n3631 0.00735484
R14672 dvss.n3633 dvss 0.00735484
R14673 dvss.n3632 dvss 0.00735484
R14674 dvss dvss.n3641 0.00735484
R14675 dvss dvss.n3642 0.00735484
R14676 dvss.n3645 dvss 0.00735484
R14677 dvss.n3644 dvss 0.00735484
R14678 dvss.n3643 dvss 0.00735484
R14679 dvss dvss.n3653 0.00735484
R14680 dvss.n3655 dvss 0.00735484
R14681 dvss.n3654 dvss 0.00735484
R14682 dvss.n3660 dvss 0.00735484
R14683 dvss.n3659 dvss 0.00735484
R14684 dvss.n493 dvss 0.00735484
R14685 dvss.n3670 dvss 0.00735484
R14686 dvss.n3669 dvss 0.00735484
R14687 dvss.n487 dvss 0.00735484
R14688 dvss.n3674 dvss 0.00735484
R14689 dvss.n484 dvss 0.00735484
R14690 dvss dvss.n3684 0.00735484
R14691 dvss dvss.n3685 0.00735484
R14692 dvss.n3686 dvss 0.00735484
R14693 dvss.n477 dvss 0.00735484
R14694 dvss.n476 dvss 0.00735484
R14695 dvss dvss.n3698 0.00735484
R14696 dvss dvss.n3699 0.00735484
R14697 dvss.n3805 dvss 0.00735484
R14698 dvss.n3804 dvss 0.00735484
R14699 dvss.n3803 dvss 0.00735484
R14700 dvss.n3800 dvss 0.00735484
R14701 dvss.n3799 dvss 0.00735484
R14702 dvss.n3798 dvss 0.00735484
R14703 dvss.n3795 dvss 0.00735484
R14704 dvss.n3794 dvss 0.00735484
R14705 dvss.n3793 dvss 0.00735484
R14706 dvss.n3707 dvss 0.00735484
R14707 dvss.n3790 dvss 0.00735484
R14708 dvss.n3789 dvss 0.00735484
R14709 dvss.n3786 dvss 0.00735484
R14710 dvss.n3785 dvss 0.00735484
R14711 dvss dvss.n3714 0.00735484
R14712 dvss.n3781 dvss 0.00735484
R14713 dvss.n3780 dvss 0.00735484
R14714 dvss.n3777 dvss 0.00735484
R14715 dvss.n3773 dvss 0.00735484
R14716 dvss.n3772 dvss 0.00735484
R14717 dvss.n3769 dvss 0.00735484
R14718 dvss.n3768 dvss 0.00735484
R14719 dvss.n3767 dvss 0.00735484
R14720 dvss.n3763 dvss 0.00735484
R14721 dvss.n3762 dvss 0.00735484
R14722 dvss.n3759 dvss 0.00735484
R14723 dvss.n3758 dvss 0.00735484
R14724 dvss.n3757 dvss 0.00735484
R14725 dvss.n4050 dvss 0.00735484
R14726 dvss.n4049 dvss 0.00735484
R14727 dvss.n4048 dvss 0.00735484
R14728 dvss.n4133 dvss.n258 0.00725676
R14729 dvss.n1077 dvss 0.00695161
R14730 dvss.n1141 dvss 0.00695161
R14731 dvss.n1542 dvss 0.00695161
R14732 dvss dvss.n1585 0.00695161
R14733 dvss.n2017 dvss 0.00695161
R14734 dvss dvss.n2060 0.00695161
R14735 dvss dvss.n2091 0.00695161
R14736 dvss dvss.n2122 0.00695161
R14737 dvss.n3675 dvss 0.00695161
R14738 dvss dvss.n3734 0.00695161
R14739 dvss.n1086 dvss.n1079 0.00654839
R14740 dvss dvss.n986 0.0064691
R14741 dvss.n948 dvss 0.0064691
R14742 dvss dvss.n1238 0.0064691
R14743 dvss.n1239 dvss 0.0064691
R14744 dvss.n1244 dvss 0.0064691
R14745 dvss.n1252 dvss 0.0064691
R14746 dvss.n1251 dvss 0.0064691
R14747 dvss dvss.n1256 0.0064691
R14748 dvss.n1257 dvss 0.0064691
R14749 dvss dvss.n1264 0.0064691
R14750 dvss.n1265 dvss 0.0064691
R14751 dvss.n1272 dvss 0.0064691
R14752 dvss.n1271 dvss 0.0064691
R14753 dvss.n1276 dvss 0.0064691
R14754 dvss.n1275 dvss 0.0064691
R14755 dvss.n1293 dvss 0.0064691
R14756 dvss.n1292 dvss 0.0064691
R14757 dvss.n1303 dvss 0.0064691
R14758 dvss.n1302 dvss 0.0064691
R14759 dvss.n1301 dvss 0.0064691
R14760 dvss.n1317 dvss 0.0064691
R14761 dvss.n1316 dvss 0.0064691
R14762 dvss.n1326 dvss 0.0064691
R14763 dvss.n1325 dvss 0.0064691
R14764 dvss.n1484 dvss 0.0064691
R14765 dvss.n1483 dvss 0.0064691
R14766 dvss.n1482 dvss 0.0064691
R14767 dvss.n1479 dvss 0.0064691
R14768 dvss.n1478 dvss 0.0064691
R14769 dvss.n1477 dvss 0.0064691
R14770 dvss.n1474 dvss 0.0064691
R14771 dvss.n1346 dvss 0.0064691
R14772 dvss.n1471 dvss 0.0064691
R14773 dvss.n1470 dvss 0.0064691
R14774 dvss dvss.n1409 0.0064691
R14775 dvss.n1410 dvss 0.0064691
R14776 dvss.n1466 dvss 0.0064691
R14777 dvss.n1465 dvss 0.0064691
R14778 dvss.n1456 dvss 0.0064691
R14779 dvss.n1462 dvss 0.0064691
R14780 dvss.n1461 dvss 0.0064691
R14781 dvss.n1454 dvss 0.0064691
R14782 dvss dvss.n1367 0.0064691
R14783 dvss.n1451 dvss 0.0064691
R14784 dvss.n1450 dvss 0.0064691
R14785 dvss.n1449 dvss 0.0064691
R14786 dvss.n1440 dvss 0.0064691
R14787 dvss.n1437 dvss 0.0064691
R14788 dvss dvss.n1679 0.0064691
R14789 dvss.n1680 dvss 0.0064691
R14790 dvss.n1704 dvss 0.0064691
R14791 dvss.n1701 dvss 0.0064691
R14792 dvss.n1700 dvss 0.0064691
R14793 dvss.n1699 dvss 0.0064691
R14794 dvss dvss.n1713 0.0064691
R14795 dvss.n1714 dvss 0.0064691
R14796 dvss.n1719 dvss 0.0064691
R14797 dvss.n1727 dvss 0.0064691
R14798 dvss.n1726 dvss 0.0064691
R14799 dvss dvss.n1731 0.0064691
R14800 dvss.n1732 dvss 0.0064691
R14801 dvss dvss.n1739 0.0064691
R14802 dvss.n1740 dvss 0.0064691
R14803 dvss.n1747 dvss 0.0064691
R14804 dvss.n1746 dvss 0.0064691
R14805 dvss.n1751 dvss 0.0064691
R14806 dvss.n1750 dvss 0.0064691
R14807 dvss.n1768 dvss 0.0064691
R14808 dvss.n1767 dvss 0.0064691
R14809 dvss.n1778 dvss 0.0064691
R14810 dvss.n1777 dvss 0.0064691
R14811 dvss.n1776 dvss 0.0064691
R14812 dvss.n1792 dvss 0.0064691
R14813 dvss.n1791 dvss 0.0064691
R14814 dvss.n1801 dvss 0.0064691
R14815 dvss.n1800 dvss 0.0064691
R14816 dvss.n1959 dvss 0.0064691
R14817 dvss.n1958 dvss 0.0064691
R14818 dvss.n1957 dvss 0.0064691
R14819 dvss.n1954 dvss 0.0064691
R14820 dvss.n1953 dvss 0.0064691
R14821 dvss.n1952 dvss 0.0064691
R14822 dvss.n1949 dvss 0.0064691
R14823 dvss.n1821 dvss 0.0064691
R14824 dvss.n1946 dvss 0.0064691
R14825 dvss.n1945 dvss 0.0064691
R14826 dvss dvss.n1884 0.0064691
R14827 dvss.n1885 dvss 0.0064691
R14828 dvss.n1941 dvss 0.0064691
R14829 dvss.n1940 dvss 0.0064691
R14830 dvss.n1931 dvss 0.0064691
R14831 dvss.n1937 dvss 0.0064691
R14832 dvss.n1936 dvss 0.0064691
R14833 dvss.n1929 dvss 0.0064691
R14834 dvss dvss.n1842 0.0064691
R14835 dvss.n1926 dvss 0.0064691
R14836 dvss.n1925 dvss 0.0064691
R14837 dvss.n1924 dvss 0.0064691
R14838 dvss.n1915 dvss 0.0064691
R14839 dvss.n1912 dvss 0.0064691
R14840 dvss dvss.n3157 0.0064691
R14841 dvss.n3158 dvss 0.0064691
R14842 dvss.n3182 dvss 0.0064691
R14843 dvss.n3179 dvss 0.0064691
R14844 dvss.n3178 dvss 0.0064691
R14845 dvss.n3177 dvss 0.0064691
R14846 dvss dvss.n3191 0.0064691
R14847 dvss.n3192 dvss 0.0064691
R14848 dvss.n3197 dvss 0.0064691
R14849 dvss.n3205 dvss 0.0064691
R14850 dvss.n3204 dvss 0.0064691
R14851 dvss dvss.n3209 0.0064691
R14852 dvss.n3210 dvss 0.0064691
R14853 dvss dvss.n3217 0.0064691
R14854 dvss.n3218 dvss 0.0064691
R14855 dvss.n3225 dvss 0.0064691
R14856 dvss.n3224 dvss 0.0064691
R14857 dvss.n3229 dvss 0.0064691
R14858 dvss.n3228 dvss 0.0064691
R14859 dvss.n3246 dvss 0.0064691
R14860 dvss.n3245 dvss 0.0064691
R14861 dvss.n3256 dvss 0.0064691
R14862 dvss.n3255 dvss 0.0064691
R14863 dvss.n3254 dvss 0.0064691
R14864 dvss.n3271 dvss 0.0064691
R14865 dvss.n3270 dvss 0.0064691
R14866 dvss.n3280 dvss 0.0064691
R14867 dvss.n3279 dvss 0.0064691
R14868 dvss.n642 dvss 0.0064691
R14869 dvss.n3302 dvss 0.0064691
R14870 dvss.n3299 dvss 0.0064691
R14871 dvss.n3298 dvss 0.0064691
R14872 dvss dvss.n3310 0.0064691
R14873 dvss.n3311 dvss 0.0064691
R14874 dvss.n3319 dvss 0.0064691
R14875 dvss.n625 dvss 0.0064691
R14876 dvss.n624 dvss 0.0064691
R14877 dvss.n3331 dvss 0.0064691
R14878 dvss.n3330 dvss 0.0064691
R14879 dvss.n3342 dvss 0.0064691
R14880 dvss.n3341 dvss 0.0064691
R14881 dvss.n3345 dvss 0.0064691
R14882 dvss.n3337 dvss 0.0064691
R14883 dvss.n3336 dvss 0.0064691
R14884 dvss.n3354 dvss 0.0064691
R14885 dvss.n3362 dvss 0.0064691
R14886 dvss.n3361 dvss 0.0064691
R14887 dvss dvss.n3369 0.0064691
R14888 dvss.n3376 dvss 0.0064691
R14889 dvss.n3375 dvss 0.0064691
R14890 dvss.n3388 dvss 0.0064691
R14891 dvss.n3387 dvss 0.0064691
R14892 dvss.n3397 dvss 0.0064691
R14893 dvss.n3396 dvss 0.0064691
R14894 dvss.n3400 dvss 0.0064691
R14895 dvss.n3415 dvss 0.0064691
R14896 dvss.n3414 dvss 0.0064691
R14897 dvss.n3413 dvss 0.0064691
R14898 dvss dvss.n3423 0.0064691
R14899 dvss.n3424 dvss 0.0064691
R14900 dvss.n3438 dvss 0.0064691
R14901 dvss.n3437 dvss 0.0064691
R14902 dvss dvss.n3433 0.0064691
R14903 dvss.n3434 dvss 0.0064691
R14904 dvss dvss.n3448 0.0064691
R14905 dvss dvss.n3449 0.0064691
R14906 dvss.n3450 dvss 0.0064691
R14907 dvss.n3461 dvss 0.0064691
R14908 dvss dvss.n3456 0.0064691
R14909 dvss.n3458 dvss 0.0064691
R14910 dvss.n3457 dvss 0.0064691
R14911 dvss.n3478 dvss 0.0064691
R14912 dvss.n3477 dvss 0.0064691
R14913 dvss.n3488 dvss 0.0064691
R14914 dvss.n3487 dvss 0.0064691
R14915 dvss.n3486 dvss 0.0064691
R14916 dvss.n3502 dvss 0.0064691
R14917 dvss.n3501 dvss 0.0064691
R14918 dvss.n3511 dvss 0.0064691
R14919 dvss.n3510 dvss 0.0064691
R14920 dvss.n3617 dvss 0.0064691
R14921 dvss.n3616 dvss 0.0064691
R14922 dvss.n3615 dvss 0.0064691
R14923 dvss.n3612 dvss 0.0064691
R14924 dvss.n3611 dvss 0.0064691
R14925 dvss.n3610 dvss 0.0064691
R14926 dvss.n3607 dvss 0.0064691
R14927 dvss.n3531 dvss 0.0064691
R14928 dvss.n3604 dvss 0.0064691
R14929 dvss.n3603 dvss 0.0064691
R14930 dvss dvss.n3549 0.0064691
R14931 dvss.n3550 dvss 0.0064691
R14932 dvss.n3599 dvss 0.0064691
R14933 dvss.n3598 dvss 0.0064691
R14934 dvss.n3589 dvss 0.0064691
R14935 dvss.n3595 dvss 0.0064691
R14936 dvss.n3594 dvss 0.0064691
R14937 dvss.n3892 dvss 0.0064691
R14938 dvss.n384 dvss 0.0064691
R14939 dvss.n3889 dvss 0.0064691
R14940 dvss.n3888 dvss 0.0064691
R14941 dvss.n3887 dvss 0.0064691
R14942 dvss.n453 dvss 0.0064691
R14943 dvss dvss.n460 0.0064691
R14944 dvss.n461 dvss 0.0064691
R14945 dvss dvss.n387 0.0064691
R14946 dvss.n3873 dvss 0.0064691
R14947 dvss.n3872 dvss 0.0064691
R14948 dvss.n3871 dvss 0.0064691
R14949 dvss.n3868 dvss 0.0064691
R14950 dvss.n3867 dvss 0.0064691
R14951 dvss.n3866 dvss 0.0064691
R14952 dvss.n3863 dvss 0.0064691
R14953 dvss.n410 dvss 0.0064691
R14954 dvss.n3860 dvss 0.0064691
R14955 dvss.n3859 dvss 0.0064691
R14956 dvss dvss.n3827 0.0064691
R14957 dvss.n3828 dvss 0.0064691
R14958 dvss.n3855 dvss 0.0064691
R14959 dvss.n3854 dvss 0.0064691
R14960 dvss.n3845 dvss 0.0064691
R14961 dvss.n3851 dvss 0.0064691
R14962 dvss.n3850 dvss 0.0064691
R14963 dvss dvss.n3935 0.0064691
R14964 dvss dvss.n3936 0.0064691
R14965 dvss.n3937 dvss 0.0064691
R14966 dvss dvss.n3946 0.0064691
R14967 dvss.n3947 dvss 0.0064691
R14968 dvss.n3953 dvss 0.0064691
R14969 dvss.n3963 dvss 0.0064691
R14970 dvss.n3962 dvss 0.0064691
R14971 dvss.n3961 dvss 0.0064691
R14972 dvss dvss.n3977 0.0064691
R14973 dvss.n3978 dvss 0.0064691
R14974 dvss dvss.n3985 0.0064691
R14975 dvss.n2849 dvss.n2426 0.00641216
R14976 dvss.n2802 dvss.n2459 0.00641216
R14977 dvss.n2755 dvss.n2495 0.00641216
R14978 dvss.n2708 dvss.n2531 0.00641216
R14979 dvss.n2661 dvss.n2567 0.00641216
R14980 dvss.n2614 dvss.n2603 0.00641216
R14981 dvss.n2956 dvss.n2298 0.00641216
R14982 dvss.n2272 dvss.n2271 0.00641216
R14983 dvss.n4099 dvss.n281 0.00641216
R14984 dvss dvss.n914 0.00611798
R14985 dvss dvss.n915 0.00611798
R14986 dvss dvss.n916 0.00611798
R14987 dvss dvss.n971 0.00611798
R14988 dvss dvss.n919 0.00611798
R14989 dvss dvss.n920 0.00611798
R14990 dvss dvss.n921 0.00611798
R14991 dvss.n987 dvss 0.00611798
R14992 dvss dvss.n924 0.00611798
R14993 dvss dvss.n925 0.00611798
R14994 dvss dvss.n929 0.00611798
R14995 dvss dvss.n930 0.00611798
R14996 dvss.n1025 dvss 0.00611798
R14997 dvss dvss.n933 0.00611798
R14998 dvss.n1029 dvss 0.00611798
R14999 dvss.n1019 dvss 0.00611798
R15000 dvss dvss.n934 0.00611798
R15001 dvss dvss.n947 0.00611798
R15002 dvss.n1288 dvss 0.00611798
R15003 dvss dvss.n1358 0.00611798
R15004 dvss.n1763 dvss 0.00611798
R15005 dvss dvss.n1833 0.00611798
R15006 dvss.n3241 dvss 0.00611798
R15007 dvss.n3357 dvss 0.00611798
R15008 dvss.n3473 dvss 0.00611798
R15009 dvss dvss.n3586 0.00611798
R15010 dvss dvss.n3842 0.00611798
R15011 dvss.n1152 dvss 0.00574194
R15012 dvss.n1553 dvss 0.00574194
R15013 dvss dvss.n1632 0.00574194
R15014 dvss.n2028 dvss 0.00574194
R15015 dvss dvss.n3110 0.00574194
R15016 dvss dvss.n3060 0.00574194
R15017 dvss dvss.n3010 0.00574194
R15018 dvss.n3686 dvss 0.00574194
R15019 dvss dvss.n3767 0.00574194
R15020 dvss dvss.n2870 0.00556757
R15021 dvss.n1001 dvss.n926 0.00541573
R15022 dvss.n1239 dvss 0.00541573
R15023 dvss dvss.n1291 0.00541573
R15024 dvss dvss.n1477 0.00541573
R15025 dvss.n1455 dvss 0.00541573
R15026 dvss.n1714 dvss 0.00541573
R15027 dvss dvss.n1766 0.00541573
R15028 dvss dvss.n1952 0.00541573
R15029 dvss.n1930 dvss 0.00541573
R15030 dvss.n3192 dvss 0.00541573
R15031 dvss dvss.n3244 0.00541573
R15032 dvss.n3311 dvss 0.00541573
R15033 dvss dvss.n3360 0.00541573
R15034 dvss.n3424 dvss 0.00541573
R15035 dvss dvss.n3476 0.00541573
R15036 dvss dvss.n3610 0.00541573
R15037 dvss.n3588 dvss 0.00541573
R15038 dvss dvss.n3866 0.00541573
R15039 dvss.n3844 dvss 0.00541573
R15040 dvss dvss.n1301 0.00506461
R15041 dvss.n1487 dvss 0.00506461
R15042 dvss dvss.n1449 0.00506461
R15043 dvss.n1683 dvss 0.00506461
R15044 dvss dvss.n1776 0.00506461
R15045 dvss.n1962 dvss 0.00506461
R15046 dvss dvss.n1924 0.00506461
R15047 dvss.n3161 dvss 0.00506461
R15048 dvss dvss.n3254 0.00506461
R15049 dvss.n3283 dvss 0.00506461
R15050 dvss dvss.n3375 0.00506461
R15051 dvss.n3401 dvss 0.00506461
R15052 dvss dvss.n3486 0.00506461
R15053 dvss.n3620 dvss 0.00506461
R15054 dvss dvss.n3887 0.00506461
R15055 dvss.n3876 dvss 0.00506461
R15056 dvss.n3947 dvss 0.00506461
R15057 dvss.n3974 dvss 0.00506461
R15058 dvss.n1155 dvss 0.00493548
R15059 dvss.n1556 dvss 0.00493548
R15060 dvss.n1629 dvss 0.00493548
R15061 dvss.n2031 dvss 0.00493548
R15062 dvss.n3107 dvss 0.00493548
R15063 dvss.n3057 dvss 0.00493548
R15064 dvss.n3007 dvss 0.00493548
R15065 dvss.n3689 dvss 0.00493548
R15066 dvss.n3764 dvss 0.00493548
R15067 dvss.n1074 dvss.n1073 0.00412903
R15068 dvss.n1089 dvss.n1088 0.00412903
R15069 dvss dvss.n1243 0.00401124
R15070 dvss.n1296 dvss.n865 0.00401124
R15071 dvss.n1475 dvss 0.00401124
R15072 dvss.n1445 dvss.n1441 0.00401124
R15073 dvss dvss.n1718 0.00401124
R15074 dvss.n1771 dvss.n756 0.00401124
R15075 dvss.n1950 dvss 0.00401124
R15076 dvss.n1920 dvss.n1916 0.00401124
R15077 dvss dvss.n3196 0.00401124
R15078 dvss.n3249 dvss.n647 0.00401124
R15079 dvss.n3315 dvss 0.00401124
R15080 dvss.n3370 dvss.n584 0.00401124
R15081 dvss.n3428 dvss 0.00401124
R15082 dvss.n3481 dvss.n521 0.00401124
R15083 dvss.n3608 dvss 0.00401124
R15084 dvss.n3883 dvss.n383 0.00401124
R15085 dvss.n3864 dvss 0.00401124
R15086 dvss.n3952 dvss.n336 0.00401124
R15087 dvss.n2826 dvss.n2445 0.00387838
R15088 dvss.n2815 dvss.n2814 0.00387838
R15089 dvss.n2779 dvss.n2481 0.00387838
R15090 dvss.n2768 dvss.n2767 0.00387838
R15091 dvss.n2732 dvss.n2517 0.00387838
R15092 dvss.n2721 dvss.n2720 0.00387838
R15093 dvss.n2685 dvss.n2553 0.00387838
R15094 dvss.n2674 dvss.n2673 0.00387838
R15095 dvss.n2638 dvss.n2589 0.00387838
R15096 dvss.n2627 dvss.n2626 0.00387838
R15097 dvss.n2923 dvss.n2922 0.00387838
R15098 dvss.n2927 dvss.n2926 0.00387838
R15099 dvss.n2230 dvss.n2229 0.00387838
R15100 dvss.n2285 dvss.n2284 0.00387838
R15101 dvss.n365 dvss.n364 0.00387838
R15102 dvss.n4112 dvss.n4111 0.00387838
R15103 dvss.n4076 dvss.n297 0.00387838
R15104 dvss.n4065 dvss.n4064 0.00387838
R15105 dvss.n1073 dvss 0.00372581
R15106 dvss dvss.n1089 0.00372581
R15107 dvss dvss.n1117 0.00372581
R15108 dvss.n1145 dvss 0.00372581
R15109 dvss dvss.n838 0.00372581
R15110 dvss dvss.n829 0.00372581
R15111 dvss.n1581 dvss 0.00372581
R15112 dvss dvss.n1637 0.00372581
R15113 dvss dvss.n729 0.00372581
R15114 dvss dvss.n720 0.00372581
R15115 dvss.n2056 dvss 0.00372581
R15116 dvss dvss.n3115 0.00372581
R15117 dvss.n2087 dvss 0.00372581
R15118 dvss dvss.n3065 0.00372581
R15119 dvss.n2118 dvss 0.00372581
R15120 dvss dvss.n3015 0.00372581
R15121 dvss dvss.n493 0.00372581
R15122 dvss dvss.n484 0.00372581
R15123 dvss.n3714 dvss 0.00372581
R15124 dvss dvss.n3772 0.00372581
R15125 dvss.n984 dvss.n983 0.00366011
R15126 dvss.n1007 dvss.n997 0.00366011
R15127 dvss.n1002 dvss 0.00330899
R15128 dvss.n1272 dvss 0.00330899
R15129 dvss.n1293 dvss 0.00330899
R15130 dvss dvss.n1465 0.00330899
R15131 dvss dvss.n1454 0.00330899
R15132 dvss.n1747 dvss 0.00330899
R15133 dvss.n1768 dvss 0.00330899
R15134 dvss dvss.n1940 0.00330899
R15135 dvss dvss.n1929 0.00330899
R15136 dvss.n3225 dvss 0.00330899
R15137 dvss.n3246 dvss 0.00330899
R15138 dvss.n3345 dvss 0.00330899
R15139 dvss.n3362 dvss 0.00330899
R15140 dvss.n3461 dvss 0.00330899
R15141 dvss.n3478 dvss 0.00330899
R15142 dvss dvss.n3598 0.00330899
R15143 dvss.n3892 dvss 0.00330899
R15144 dvss dvss.n3854 0.00330899
R15145 dvss.n3935 dvss 0.00330899
R15146 dvss dvss.n2817 0.00303378
R15147 dvss dvss.n2770 0.00303378
R15148 dvss dvss.n2723 0.00303378
R15149 dvss dvss.n2676 0.00303378
R15150 dvss dvss.n2629 0.00303378
R15151 dvss dvss.n2929 0.00303378
R15152 dvss dvss.n2216 0.00303378
R15153 dvss dvss.n271 0.00303378
R15154 dvss dvss.n4067 0.00303378
R15155 dvss.n982 dvss 0.00295787
R15156 dvss dvss.n1008 0.00295787
R15157 dvss.n1243 dvss.n901 0.00295787
R15158 dvss.n868 dvss 0.00295787
R15159 dvss.n1296 dvss 0.00295787
R15160 dvss.n1475 dvss.n1339 0.00295787
R15161 dvss.n1446 dvss 0.00295787
R15162 dvss.n1441 dvss 0.00295787
R15163 dvss.n1718 dvss.n792 0.00295787
R15164 dvss.n759 dvss 0.00295787
R15165 dvss.n1771 dvss 0.00295787
R15166 dvss.n1950 dvss.n1814 0.00295787
R15167 dvss.n1921 dvss 0.00295787
R15168 dvss.n1916 dvss 0.00295787
R15169 dvss.n3196 dvss.n683 0.00295787
R15170 dvss.n650 dvss 0.00295787
R15171 dvss.n3249 dvss 0.00295787
R15172 dvss.n3316 dvss.n3315 0.00295787
R15173 dvss.n587 dvss 0.00295787
R15174 dvss.n3370 dvss 0.00295787
R15175 dvss.n3429 dvss.n3428 0.00295787
R15176 dvss.n524 dvss 0.00295787
R15177 dvss.n3481 dvss 0.00295787
R15178 dvss.n3608 dvss.n3524 0.00295787
R15179 dvss.n3884 dvss 0.00295787
R15180 dvss dvss.n383 0.00295787
R15181 dvss.n3864 dvss.n403 0.00295787
R15182 dvss.n339 dvss 0.00295787
R15183 dvss dvss.n3952 0.00295787
R15184 dvss.n1130 dvss 0.00291935
R15185 dvss.n1155 dvss.n1154 0.00291935
R15186 dvss.n1522 dvss 0.00291935
R15187 dvss.n1557 dvss.n1556 0.00291935
R15188 dvss.n1655 dvss 0.00291935
R15189 dvss.n1629 dvss.n1591 0.00291935
R15190 dvss.n1997 dvss 0.00291935
R15191 dvss.n2032 dvss.n2031 0.00291935
R15192 dvss.n3133 dvss 0.00291935
R15193 dvss.n3107 dvss.n2066 0.00291935
R15194 dvss.n3083 dvss 0.00291935
R15195 dvss.n3057 dvss.n2097 0.00291935
R15196 dvss.n3033 dvss 0.00291935
R15197 dvss.n3007 dvss.n2128 0.00291935
R15198 dvss.n3655 dvss 0.00291935
R15199 dvss.n3690 dvss.n3689 0.00291935
R15200 dvss.n3790 dvss 0.00291935
R15201 dvss.n3764 dvss.n3740 0.00291935
R15202 dvss.n1002 dvss 0.00260674
R15203 dvss.n1256 dvss 0.00260674
R15204 dvss.n1320 dvss.n868 0.00260674
R15205 dvss dvss.n1470 0.00260674
R15206 dvss.n1446 dvss.n1372 0.00260674
R15207 dvss.n1731 dvss 0.00260674
R15208 dvss.n1795 dvss.n759 0.00260674
R15209 dvss dvss.n1945 0.00260674
R15210 dvss.n1921 dvss.n1847 0.00260674
R15211 dvss.n3209 dvss 0.00260674
R15212 dvss.n3274 dvss.n650 0.00260674
R15213 dvss.n3331 dvss 0.00260674
R15214 dvss.n3391 dvss.n587 0.00260674
R15215 dvss.n3434 dvss 0.00260674
R15216 dvss.n3505 dvss.n524 0.00260674
R15217 dvss dvss.n3603 0.00260674
R15218 dvss.n3884 dvss.n382 0.00260674
R15219 dvss dvss.n3859 0.00260674
R15220 dvss.n3956 dvss.n339 0.00260674
R15221 dvss.n1321 dvss.n1320 0.00190449
R15222 dvss.n1487 dvss.n860 0.00190449
R15223 dvss.n1443 dvss.n1372 0.00190449
R15224 dvss.n1683 dvss.n1682 0.00190449
R15225 dvss.n1796 dvss.n1795 0.00190449
R15226 dvss.n1962 dvss.n751 0.00190449
R15227 dvss.n1918 dvss.n1847 0.00190449
R15228 dvss.n3161 dvss.n3160 0.00190449
R15229 dvss.n3275 dvss.n3274 0.00190449
R15230 dvss.n3283 dvss.n641 0.00190449
R15231 dvss.n3392 dvss.n3391 0.00190449
R15232 dvss.n3401 dvss.n579 0.00190449
R15233 dvss.n3506 dvss.n3505 0.00190449
R15234 dvss.n3620 dvss.n516 0.00190449
R15235 dvss.n3881 dvss.n382 0.00190449
R15236 dvss.n3877 dvss.n3876 0.00190449
R15237 dvss.n3957 dvss.n3956 0.00190449
R15238 dvss.n3974 dvss.n322 0.00190449
R15239 dvss.n1291 dvss.n881 0.00155337
R15240 dvss dvss.n1325 0.00155337
R15241 dvss.n1455 dvss.n1359 0.00155337
R15242 dvss.n1680 dvss 0.00155337
R15243 dvss.n1766 dvss.n772 0.00155337
R15244 dvss dvss.n1800 0.00155337
R15245 dvss.n1930 dvss.n1834 0.00155337
R15246 dvss.n3158 dvss 0.00155337
R15247 dvss.n3244 dvss.n663 0.00155337
R15248 dvss dvss.n3279 0.00155337
R15249 dvss.n3360 dvss.n603 0.00155337
R15250 dvss dvss.n3396 0.00155337
R15251 dvss.n3476 dvss.n537 0.00155337
R15252 dvss dvss.n3510 0.00155337
R15253 dvss.n3588 dvss.n3587 0.00155337
R15254 dvss dvss.n387 0.00155337
R15255 dvss.n3844 dvss.n3843 0.00155337
R15256 dvss dvss.n3961 0.00155337
R15257 dvss.n2868 dvss.n2867 0.00134459
R15258 dvss.n1086 dvss 0.00130645
R15259 dvss dvss.n1001 0.00120225
R15260 dvss.n1142 dvss.n1141 0.000903226
R15261 dvss.n1160 dvss 0.000903226
R15262 dvss.n1542 dvss.n828 0.000903226
R15263 dvss dvss.n821 0.000903226
R15264 dvss.n1641 dvss.n1585 0.000903226
R15265 dvss dvss.n1627 0.000903226
R15266 dvss.n2017 dvss.n719 0.000903226
R15267 dvss dvss.n712 0.000903226
R15268 dvss.n3119 dvss.n2060 0.000903226
R15269 dvss dvss.n3105 0.000903226
R15270 dvss.n3069 dvss.n2091 0.000903226
R15271 dvss dvss.n3055 0.000903226
R15272 dvss.n3019 dvss.n2122 0.000903226
R15273 dvss dvss.n3005 0.000903226
R15274 dvss.n3675 dvss.n483 0.000903226
R15275 dvss dvss.n476 0.000903226
R15276 dvss.n3776 dvss.n3734 0.000903226
R15277 dvss dvss.n3762 0.000903226
R15278 dvss.n961 dvss.n915 0.000851124
R15279 dvss.n959 dvss.n916 0.000851124
R15280 dvss.n971 dvss.n970 0.000851124
R15281 dvss.n972 dvss.n919 0.000851124
R15282 dvss.n974 dvss.n920 0.000851124
R15283 dvss.n956 dvss.n921 0.000851124
R15284 dvss.n983 dvss.n982 0.000851124
R15285 dvss.n987 dvss.n924 0.000851124
R15286 dvss.n989 dvss.n925 0.000851124
R15287 dvss.n953 dvss.n926 0.000851124
R15288 dvss.n1008 dvss.n1007 0.000851124
R15289 dvss.n1009 dvss.n929 0.000851124
R15290 dvss.n1011 dvss.n930 0.000851124
R15291 dvss.n1026 dvss.n1025 0.000851124
R15292 dvss.n1029 dvss.n933 0.000851124
R15293 dvss.n1028 dvss.n1019 0.000851124
R15294 dvss.n1018 dvss.n934 0.000851124
R15295 dvss.n947 dvss.n939 0.000851124
R15296 dvss.n1289 dvss.n1288 0.000851124
R15297 dvss.n1317 dvss 0.000851124
R15298 dvss.n1460 dvss.n1358 0.000851124
R15299 dvss dvss.n1440 0.000851124
R15300 dvss.n1764 dvss.n1763 0.000851124
R15301 dvss.n1792 dvss 0.000851124
R15302 dvss.n1935 dvss.n1833 0.000851124
R15303 dvss dvss.n1915 0.000851124
R15304 dvss.n3242 dvss.n3241 0.000851124
R15305 dvss.n3271 dvss 0.000851124
R15306 dvss.n3358 dvss.n3357 0.000851124
R15307 dvss.n3388 dvss 0.000851124
R15308 dvss.n3474 dvss.n3473 0.000851124
R15309 dvss.n3502 dvss 0.000851124
R15310 dvss.n3593 dvss.n3586 0.000851124
R15311 dvss.n453 dvss 0.000851124
R15312 dvss.n3849 dvss.n3842 0.000851124
R15313 dvss.n3953 dvss 0.000851124
R15314 rc_osc_0.n.n4 rc_osc_0.n.t6 244.843
R15315 rc_osc_0.n.n2 rc_osc_0.n.t11 240.778
R15316 rc_osc_0.n.n3 rc_osc_0.n.t13 240.349
R15317 rc_osc_0.n.n2 rc_osc_0.n.t9 240.349
R15318 rc_osc_0.n.n10 rc_osc_0.n.n0 211.296
R15319 rc_osc_0.n.n11 rc_osc_0.n.n10 204.284
R15320 rc_osc_0.n.n7 rc_osc_0.n.t10 123.462
R15321 rc_osc_0.n.n5 rc_osc_0.n.t7 120.871
R15322 rc_osc_0.n.n6 rc_osc_0.n.t8 120.773
R15323 rc_osc_0.n.n5 rc_osc_0.n.t12 120.174
R15324 rc_osc_0.n.n9 rc_osc_0.n.n1 72.3553
R15325 rc_osc_0.n.n0 rc_osc_0.n.t1 28.5655
R15326 rc_osc_0.n.n0 rc_osc_0.n.t2 28.5655
R15327 rc_osc_0.n.n11 rc_osc_0.n.t3 28.5655
R15328 rc_osc_0.n.t0 rc_osc_0.n.n11 28.5655
R15329 rc_osc_0.n.n1 rc_osc_0.n.t5 17.4005
R15330 rc_osc_0.n.n1 rc_osc_0.n.t4 17.4005
R15331 rc_osc_0.n.n4 rc_osc_0.n.n3 9.0153
R15332 rc_osc_0.n.n7 rc_osc_0.n.n6 5.23012
R15333 rc_osc_0.n.n8 rc_osc_0.n.n7 3.78258
R15334 rc_osc_0.n.n9 rc_osc_0.n.n8 3.4105
R15335 rc_osc_0.n.n10 rc_osc_0.n.n9 1.35184
R15336 rc_osc_0.n.n3 rc_osc_0.n.n2 0.408448
R15337 rc_osc_0.n.n8 rc_osc_0.n.n4 0.147461
R15338 rc_osc_0.n.n6 rc_osc_0.n.n5 0.049413
R15339 brout_filt.n2 brout_filt.n0 243.458
R15340 brout_filt.n2 brout_filt.n1 205.059
R15341 brout_filt.n4 brout_filt.n3 205.059
R15342 brout_filt.n6 brout_filt.n5 205.059
R15343 brout_filt.n8 brout_filt.n7 205.059
R15344 brout_filt.n10 brout_filt.n9 205.059
R15345 brout_filt.n12 brout_filt.n11 205.059
R15346 brout_filt.n14 brout_filt.n13 205.059
R15347 brout_filt.n18 brout_filt.n16 133.534
R15348 brout_filt.n18 brout_filt.n17 99.1759
R15349 brout_filt.n20 brout_filt.n19 99.1759
R15350 brout_filt.n22 brout_filt.n21 99.1759
R15351 brout_filt.n24 brout_filt.n23 99.1759
R15352 brout_filt.n26 brout_filt.n25 99.1759
R15353 brout_filt.n28 brout_filt.n27 99.1759
R15354 brout_filt brout_filt.n29 97.4305
R15355 brout_filt.n4 brout_filt.n2 38.4005
R15356 brout_filt.n6 brout_filt.n4 38.4005
R15357 brout_filt.n8 brout_filt.n6 38.4005
R15358 brout_filt.n10 brout_filt.n8 38.4005
R15359 brout_filt.n12 brout_filt.n10 38.4005
R15360 brout_filt.n14 brout_filt.n12 38.4005
R15361 brout_filt.n20 brout_filt.n18 34.3584
R15362 brout_filt.n22 brout_filt.n20 34.3584
R15363 brout_filt.n24 brout_filt.n22 34.3584
R15364 brout_filt.n26 brout_filt.n24 34.3584
R15365 brout_filt.n28 brout_filt.n26 34.3584
R15366 brout_filt.n30 brout_filt.n28 34.3584
R15367 brout_filt.n13 brout_filt.t3 26.5955
R15368 brout_filt.n13 brout_filt.t9 26.5955
R15369 brout_filt.n0 brout_filt.t1 26.5955
R15370 brout_filt.n0 brout_filt.t8 26.5955
R15371 brout_filt.n1 brout_filt.t15 26.5955
R15372 brout_filt.n1 brout_filt.t11 26.5955
R15373 brout_filt.n3 brout_filt.t14 26.5955
R15374 brout_filt.n3 brout_filt.t6 26.5955
R15375 brout_filt.n5 brout_filt.t2 26.5955
R15376 brout_filt.n5 brout_filt.t5 26.5955
R15377 brout_filt.n7 brout_filt.t13 26.5955
R15378 brout_filt.n7 brout_filt.t7 26.5955
R15379 brout_filt.n9 brout_filt.t0 26.5955
R15380 brout_filt.n9 brout_filt.t12 26.5955
R15381 brout_filt.n11 brout_filt.t4 26.5955
R15382 brout_filt.n11 brout_filt.t10 26.5955
R15383 brout_filt.n29 brout_filt.t30 24.9236
R15384 brout_filt.n29 brout_filt.t20 24.9236
R15385 brout_filt.n16 brout_filt.t28 24.9236
R15386 brout_filt.n16 brout_filt.t19 24.9236
R15387 brout_filt.n17 brout_filt.t26 24.9236
R15388 brout_filt.n17 brout_filt.t22 24.9236
R15389 brout_filt.n19 brout_filt.t25 24.9236
R15390 brout_filt.n19 brout_filt.t17 24.9236
R15391 brout_filt.n21 brout_filt.t29 24.9236
R15392 brout_filt.n21 brout_filt.t16 24.9236
R15393 brout_filt.n23 brout_filt.t24 24.9236
R15394 brout_filt.n23 brout_filt.t18 24.9236
R15395 brout_filt.n25 brout_filt.t27 24.9236
R15396 brout_filt.n25 brout_filt.t23 24.9236
R15397 brout_filt.n27 brout_filt.t31 24.9236
R15398 brout_filt.n27 brout_filt.t21 24.9236
R15399 brout_filt.n15 brout_filt.n14 12.6066
R15400 brout_filt brout_filt.n30 11.4429
R15401 brout_filt brout_filt.n15 5.81868
R15402 brout_filt.n15 brout_filt 4.52868
R15403 brout_filt.n30 brout_filt 1.74595
R15404 rstring_mux_0.vtop.n4 rstring_mux_0.vtop.t0 87.3599
R15405 rstring_mux_0.vtop.n2 rstring_mux_0.vtop.n0 48.5415
R15406 rstring_mux_0.vtop.n13 rstring_mux_0.vtop.n12 48.4284
R15407 rstring_mux_0.vtop.n11 rstring_mux_0.vtop.n10 48.4284
R15408 rstring_mux_0.vtop.n9 rstring_mux_0.vtop.n8 48.4284
R15409 rstring_mux_0.vtop.n7 rstring_mux_0.vtop.n6 48.4284
R15410 rstring_mux_0.vtop.n2 rstring_mux_0.vtop.n1 48.4284
R15411 rstring_mux_0.vtop.n15 rstring_mux_0.vtop.n14 45.0184
R15412 rstring_mux_0.vtop.n4 rstring_mux_0.vtop.n3 45.0184
R15413 rstring_mux_0.vtop rstring_mux_0.vtop.t17 19.1879
R15414 rstring_mux_0.vtop.n14 rstring_mux_0.vtop.t4 5.5395
R15415 rstring_mux_0.vtop.n14 rstring_mux_0.vtop.t11 5.5395
R15416 rstring_mux_0.vtop.n12 rstring_mux_0.vtop.t5 5.5395
R15417 rstring_mux_0.vtop.n12 rstring_mux_0.vtop.t13 5.5395
R15418 rstring_mux_0.vtop.n10 rstring_mux_0.vtop.t7 5.5395
R15419 rstring_mux_0.vtop.n10 rstring_mux_0.vtop.t15 5.5395
R15420 rstring_mux_0.vtop.n8 rstring_mux_0.vtop.t2 5.5395
R15421 rstring_mux_0.vtop.n8 rstring_mux_0.vtop.t9 5.5395
R15422 rstring_mux_0.vtop.n6 rstring_mux_0.vtop.t3 5.5395
R15423 rstring_mux_0.vtop.n6 rstring_mux_0.vtop.t10 5.5395
R15424 rstring_mux_0.vtop.n3 rstring_mux_0.vtop.t14 5.5395
R15425 rstring_mux_0.vtop.n3 rstring_mux_0.vtop.t12 5.5395
R15426 rstring_mux_0.vtop.n1 rstring_mux_0.vtop.t16 5.5395
R15427 rstring_mux_0.vtop.n1 rstring_mux_0.vtop.t6 5.5395
R15428 rstring_mux_0.vtop.n0 rstring_mux_0.vtop.t1 5.5395
R15429 rstring_mux_0.vtop.n0 rstring_mux_0.vtop.t8 5.5395
R15430 rstring_mux_0.vtop.n15 rstring_mux_0.vtop.n13 3.5118
R15431 rstring_mux_0.vtop.n5 rstring_mux_0.vtop.n4 3.4105
R15432 rstring_mux_0.vtop rstring_mux_0.vtop.n15 0.829892
R15433 rstring_mux_0.vtop.n5 rstring_mux_0.vtop.n2 0.113554
R15434 rstring_mux_0.vtop.n7 rstring_mux_0.vtop.n5 0.113554
R15435 rstring_mux_0.vtop.n9 rstring_mux_0.vtop.n7 0.113554
R15436 rstring_mux_0.vtop.n11 rstring_mux_0.vtop.n9 0.113554
R15437 rstring_mux_0.vtop.n13 rstring_mux_0.vtop.n11 0.113554
R15438 otrip_decoded[0].n0 otrip_decoded[0].t1 186.374
R15439 otrip_decoded[0].n0 otrip_decoded[0].t0 170.308
R15440 otrip_decoded[0] otrip_decoded[0].n1 154.56
R15441 otrip_decoded[0].n2 otrip_decoded[0].n1 153.462
R15442 otrip_decoded[0].n1 otrip_decoded[0].n0 101.513
R15443 otrip_decoded[0].n3 otrip_decoded[0] 11.8005
R15444 otrip_decoded[0].n3 otrip_decoded[0].n2 4.96991
R15445 otrip_decoded[0].n2 otrip_decoded[0] 3.46403
R15446 otrip_decoded[0] otrip_decoded[0].n3 2.71109
R15447 dcomp.n2 dcomp.n0 243.458
R15448 dcomp.n2 dcomp.n1 205.059
R15449 dcomp.n4 dcomp.n3 205.059
R15450 dcomp.n6 dcomp.n5 205.059
R15451 dcomp.n8 dcomp.n7 205.059
R15452 dcomp.n10 dcomp.n9 205.059
R15453 dcomp.n12 dcomp.n11 205.059
R15454 dcomp.n14 dcomp.n13 205.059
R15455 dcomp.n17 dcomp.n15 133.534
R15456 dcomp.n17 dcomp.n16 99.1759
R15457 dcomp.n19 dcomp.n18 99.1759
R15458 dcomp.n21 dcomp.n20 99.1759
R15459 dcomp.n23 dcomp.n22 99.1759
R15460 dcomp.n25 dcomp.n24 99.1759
R15461 dcomp.n27 dcomp.n26 99.1759
R15462 dcomp dcomp.n28 97.4305
R15463 dcomp.n4 dcomp.n2 38.4005
R15464 dcomp.n6 dcomp.n4 38.4005
R15465 dcomp.n8 dcomp.n6 38.4005
R15466 dcomp.n10 dcomp.n8 38.4005
R15467 dcomp.n12 dcomp.n10 38.4005
R15468 dcomp.n14 dcomp.n12 38.4005
R15469 dcomp.n19 dcomp.n17 34.3584
R15470 dcomp.n21 dcomp.n19 34.3584
R15471 dcomp.n23 dcomp.n21 34.3584
R15472 dcomp.n25 dcomp.n23 34.3584
R15473 dcomp.n27 dcomp.n25 34.3584
R15474 dcomp.n29 dcomp.n27 34.3584
R15475 dcomp.n13 dcomp.t10 26.5955
R15476 dcomp.n13 dcomp.t0 26.5955
R15477 dcomp.n0 dcomp.t8 26.5955
R15478 dcomp.n0 dcomp.t15 26.5955
R15479 dcomp.n1 dcomp.t6 26.5955
R15480 dcomp.n1 dcomp.t2 26.5955
R15481 dcomp.n3 dcomp.t5 26.5955
R15482 dcomp.n3 dcomp.t13 26.5955
R15483 dcomp.n5 dcomp.t9 26.5955
R15484 dcomp.n5 dcomp.t12 26.5955
R15485 dcomp.n7 dcomp.t4 26.5955
R15486 dcomp.n7 dcomp.t14 26.5955
R15487 dcomp.n9 dcomp.t7 26.5955
R15488 dcomp.n9 dcomp.t3 26.5955
R15489 dcomp.n11 dcomp.t11 26.5955
R15490 dcomp.n11 dcomp.t1 26.5955
R15491 dcomp.n28 dcomp.t20 24.9236
R15492 dcomp.n28 dcomp.t26 24.9236
R15493 dcomp.n15 dcomp.t18 24.9236
R15494 dcomp.n15 dcomp.t25 24.9236
R15495 dcomp.n16 dcomp.t16 24.9236
R15496 dcomp.n16 dcomp.t28 24.9236
R15497 dcomp.n18 dcomp.t31 24.9236
R15498 dcomp.n18 dcomp.t23 24.9236
R15499 dcomp.n20 dcomp.t19 24.9236
R15500 dcomp.n20 dcomp.t22 24.9236
R15501 dcomp.n22 dcomp.t30 24.9236
R15502 dcomp.n22 dcomp.t24 24.9236
R15503 dcomp.n24 dcomp.t17 24.9236
R15504 dcomp.n24 dcomp.t29 24.9236
R15505 dcomp.n26 dcomp.t21 24.9236
R15506 dcomp.n26 dcomp.t27 24.9236
R15507 dcomp dcomp.n14 18.4247
R15508 dcomp.n30 dcomp.n29 10.0853
R15509 dcomp.n30 dcomp 4.84706
R15510 dcomp.n29 dcomp 1.74595
R15511 dcomp dcomp.n30 1.35808
R15512 schmitt_trigger_0.in.n3 schmitt_trigger_0.in.t2 240.778
R15513 schmitt_trigger_0.in.n0 schmitt_trigger_0.in.t8 240.778
R15514 schmitt_trigger_0.in.n3 schmitt_trigger_0.in.t9 240.349
R15515 schmitt_trigger_0.in.n2 schmitt_trigger_0.in.t4 240.349
R15516 schmitt_trigger_0.in.n1 schmitt_trigger_0.in.t1 240.349
R15517 schmitt_trigger_0.in.n0 schmitt_trigger_0.in.t10 240.349
R15518 schmitt_trigger_0.in.n12 schmitt_trigger_0.in.t3 236.423
R15519 schmitt_trigger_0.in.n12 schmitt_trigger_0.in.t5 236.011
R15520 schmitt_trigger_0.in.n10 schmitt_trigger_0.in.n9 28.545
R15521 schmitt_trigger_0.in.n11 schmitt_trigger_0.in.n10 19.9248
R15522 schmitt_trigger_0.in.n10 schmitt_trigger_0.in.t0 5.93425
R15523 schmitt_trigger_0.in schmitt_trigger_0.in.n12 4.93075
R15524 schmitt_trigger_0.in.n11 schmitt_trigger_0.in.n4 4.72087
R15525 schmitt_trigger_0.in.n1 schmitt_trigger_0.in.n0 0.429848
R15526 schmitt_trigger_0.in.n2 schmitt_trigger_0.in.n1 0.429848
R15527 schmitt_trigger_0.in.n4 schmitt_trigger_0.in.n2 0.285826
R15528 schmitt_trigger_0.in schmitt_trigger_0.in.n11 0.216402
R15529 schmitt_trigger_0.in.n4 schmitt_trigger_0.in.n3 0.0956087
R15530 schmitt_trigger_0.in.n5 schmitt_trigger_0.in.t7 0.0791747
R15531 schmitt_trigger_0.in.n6 schmitt_trigger_0.in.n5 0.06865
R15532 schmitt_trigger_0.in.n7 schmitt_trigger_0.in.n6 0.06865
R15533 schmitt_trigger_0.in.n8 schmitt_trigger_0.in.n7 0.06865
R15534 schmitt_trigger_0.in.n9 schmitt_trigger_0.in.n8 0.06865
R15535 schmitt_trigger_0.in.n5 schmitt_trigger_0.in.t14 0.0110247
R15536 schmitt_trigger_0.in.n6 schmitt_trigger_0.in.t12 0.0110247
R15537 schmitt_trigger_0.in.n7 schmitt_trigger_0.in.t6 0.0110247
R15538 schmitt_trigger_0.in.n8 schmitt_trigger_0.in.t13 0.0110247
R15539 schmitt_trigger_0.in.n9 schmitt_trigger_0.in.t11 0.0110247
R15540 schmitt_trigger_0.m.n5 schmitt_trigger_0.m.t15 240.764
R15541 schmitt_trigger_0.m.n6 schmitt_trigger_0.m.t16 240.713
R15542 schmitt_trigger_0.m.n7 schmitt_trigger_0.m.t17 240.529
R15543 schmitt_trigger_0.m.n5 schmitt_trigger_0.m.t14 240.349
R15544 schmitt_trigger_0.m.n10 schmitt_trigger_0.m.n8 211.214
R15545 schmitt_trigger_0.m.n2 schmitt_trigger_0.m.n0 207.804
R15546 schmitt_trigger_0.m.n2 schmitt_trigger_0.m.n1 207.585
R15547 schmitt_trigger_0.m.n4 schmitt_trigger_0.m.n3 204.175
R15548 schmitt_trigger_0.m.n10 schmitt_trigger_0.m.n9 204.175
R15549 schmitt_trigger_0.m.n13 schmitt_trigger_0.m.n12 70.9014
R15550 schmitt_trigger_0.m.n15 schmitt_trigger_0.m.n14 70.9014
R15551 schmitt_trigger_0.m.n8 schmitt_trigger_0.m.t12 28.5655
R15552 schmitt_trigger_0.m.n8 schmitt_trigger_0.m.t10 28.5655
R15553 schmitt_trigger_0.m.n3 schmitt_trigger_0.m.t1 28.5655
R15554 schmitt_trigger_0.m.n3 schmitt_trigger_0.m.t4 28.5655
R15555 schmitt_trigger_0.m.n1 schmitt_trigger_0.m.t5 28.5655
R15556 schmitt_trigger_0.m.n1 schmitt_trigger_0.m.t3 28.5655
R15557 schmitt_trigger_0.m.n0 schmitt_trigger_0.m.t2 28.5655
R15558 schmitt_trigger_0.m.n0 schmitt_trigger_0.m.t0 28.5655
R15559 schmitt_trigger_0.m.n9 schmitt_trigger_0.m.t9 28.5655
R15560 schmitt_trigger_0.m.n9 schmitt_trigger_0.m.t8 28.5655
R15561 schmitt_trigger_0.m.n12 schmitt_trigger_0.m.t13 17.4005
R15562 schmitt_trigger_0.m.n12 schmitt_trigger_0.m.t11 17.4005
R15563 schmitt_trigger_0.m.n14 schmitt_trigger_0.m.t6 17.4005
R15564 schmitt_trigger_0.m.n14 schmitt_trigger_0.m.t7 17.4005
R15565 schmitt_trigger_0.m.n7 schmitt_trigger_0.m.n6 12.9318
R15566 schmitt_trigger_0.m.n11 schmitt_trigger_0.m.n10 8.3606
R15567 schmitt_trigger_0.m.n4 schmitt_trigger_0.m.n2 3.62811
R15568 schmitt_trigger_0.m schmitt_trigger_0.m.n4 0.819515
R15569 schmitt_trigger_0.m schmitt_trigger_0.m.n15 0.73133
R15570 schmitt_trigger_0.m.n15 schmitt_trigger_0.m.n13 0.688
R15571 schmitt_trigger_0.m.n11 schmitt_trigger_0.m.n7 0.358635
R15572 schmitt_trigger_0.m.n13 schmitt_trigger_0.m.n11 0.251558
R15573 schmitt_trigger_0.m.n6 schmitt_trigger_0.m.n5 0.0297969
R15574 vbg_1v2.n68 vbg_1v2.t34 384.709
R15575 vbg_1v2.n67 vbg_1v2.t34 384.709
R15576 vbg_1v2.n78 vbg_1v2.t13 384.226
R15577 vbg_1v2.t13 vbg_1v2.n63 384.226
R15578 vbg_1v2.n77 vbg_1v2.t41 384.226
R15579 vbg_1v2.t41 vbg_1v2.n76 384.226
R15580 vbg_1v2.t3 vbg_1v2.n64 384.226
R15581 vbg_1v2.n75 vbg_1v2.t3 384.226
R15582 vbg_1v2.t5 vbg_1v2.n73 384.226
R15583 vbg_1v2.n74 vbg_1v2.t5 384.226
R15584 vbg_1v2.n72 vbg_1v2.t8 384.226
R15585 vbg_1v2.t8 vbg_1v2.n65 384.226
R15586 vbg_1v2.n71 vbg_1v2.t15 384.226
R15587 vbg_1v2.t15 vbg_1v2.n70 384.226
R15588 vbg_1v2.t20 vbg_1v2.n66 384.226
R15589 vbg_1v2.n69 vbg_1v2.t20 384.226
R15590 vbg_1v2.t30 vbg_1v2.n67 384.226
R15591 vbg_1v2.n68 vbg_1v2.t30 384.226
R15592 vbg_1v2.t22 vbg_1v2.n79 384.226
R15593 vbg_1v2.n80 vbg_1v2.t22 384.226
R15594 vbg_1v2.n62 vbg_1v2.n61 48.1045
R15595 vbg_1v2 vbg_1v2.n30 30.7468
R15596 vbg_1v2.n29 vbg_1v2.t40 14.8978
R15597 vbg_1v2.n28 vbg_1v2.t40 14.8978
R15598 vbg_1v2.n25 vbg_1v2.t25 14.8978
R15599 vbg_1v2.n24 vbg_1v2.t25 14.8978
R15600 vbg_1v2.n21 vbg_1v2.t17 14.8978
R15601 vbg_1v2.n20 vbg_1v2.t17 14.8978
R15602 vbg_1v2.n17 vbg_1v2.t1 14.8978
R15603 vbg_1v2.n16 vbg_1v2.t1 14.8978
R15604 vbg_1v2.n13 vbg_1v2.t18 14.8978
R15605 vbg_1v2.n12 vbg_1v2.t18 14.8978
R15606 vbg_1v2.n9 vbg_1v2.t2 14.8978
R15607 vbg_1v2.n8 vbg_1v2.t2 14.8978
R15608 vbg_1v2.n5 vbg_1v2.t28 14.8978
R15609 vbg_1v2.n4 vbg_1v2.t28 14.8978
R15610 vbg_1v2.n1 vbg_1v2.t21 14.8978
R15611 vbg_1v2.t21 vbg_1v2.n0 14.8978
R15612 vbg_1v2.n60 vbg_1v2.t12 14.8978
R15613 vbg_1v2.n59 vbg_1v2.t12 14.8978
R15614 vbg_1v2.n56 vbg_1v2.t14 14.8978
R15615 vbg_1v2.n55 vbg_1v2.t14 14.8978
R15616 vbg_1v2.n52 vbg_1v2.t24 14.8978
R15617 vbg_1v2.n51 vbg_1v2.t24 14.8978
R15618 vbg_1v2.n48 vbg_1v2.t4 14.8978
R15619 vbg_1v2.n47 vbg_1v2.t4 14.8978
R15620 vbg_1v2.n44 vbg_1v2.t23 14.8978
R15621 vbg_1v2.n43 vbg_1v2.t23 14.8978
R15622 vbg_1v2.n40 vbg_1v2.t36 14.8978
R15623 vbg_1v2.n39 vbg_1v2.t36 14.8978
R15624 vbg_1v2.n36 vbg_1v2.t11 14.8978
R15625 vbg_1v2.n35 vbg_1v2.t11 14.8978
R15626 vbg_1v2.n32 vbg_1v2.t19 14.8978
R15627 vbg_1v2.t19 vbg_1v2.n31 14.8978
R15628 vbg_1v2.t6 vbg_1v2.n28 12.9902
R15629 vbg_1v2.n29 vbg_1v2.t6 12.9902
R15630 vbg_1v2.t37 vbg_1v2.n24 12.9902
R15631 vbg_1v2.n25 vbg_1v2.t37 12.9902
R15632 vbg_1v2.t29 vbg_1v2.n20 12.9902
R15633 vbg_1v2.n21 vbg_1v2.t29 12.9902
R15634 vbg_1v2.t9 vbg_1v2.n16 12.9902
R15635 vbg_1v2.n17 vbg_1v2.t9 12.9902
R15636 vbg_1v2.t31 vbg_1v2.n12 12.9902
R15637 vbg_1v2.n13 vbg_1v2.t31 12.9902
R15638 vbg_1v2.t10 vbg_1v2.n8 12.9902
R15639 vbg_1v2.n9 vbg_1v2.t10 12.9902
R15640 vbg_1v2.t0 vbg_1v2.n4 12.9902
R15641 vbg_1v2.n5 vbg_1v2.t0 12.9902
R15642 vbg_1v2.t33 vbg_1v2.n0 12.9902
R15643 vbg_1v2.n1 vbg_1v2.t33 12.9902
R15644 vbg_1v2.t27 vbg_1v2.n59 12.9902
R15645 vbg_1v2.n60 vbg_1v2.t27 12.9902
R15646 vbg_1v2.t32 vbg_1v2.n55 12.9902
R15647 vbg_1v2.n56 vbg_1v2.t32 12.9902
R15648 vbg_1v2.t39 vbg_1v2.n51 12.9902
R15649 vbg_1v2.n52 vbg_1v2.t39 12.9902
R15650 vbg_1v2.t16 vbg_1v2.n47 12.9902
R15651 vbg_1v2.n48 vbg_1v2.t16 12.9902
R15652 vbg_1v2.t38 vbg_1v2.n43 12.9902
R15653 vbg_1v2.n44 vbg_1v2.t38 12.9902
R15654 vbg_1v2.t7 vbg_1v2.n39 12.9902
R15655 vbg_1v2.n40 vbg_1v2.t7 12.9902
R15656 vbg_1v2.t26 vbg_1v2.n35 12.9902
R15657 vbg_1v2.n36 vbg_1v2.t26 12.9902
R15658 vbg_1v2.t35 vbg_1v2.n31 12.9902
R15659 vbg_1v2.n32 vbg_1v2.t35 12.9902
R15660 vbg_1v2.n2 vbg_1v2.n0 5.24569
R15661 vbg_1v2.n33 vbg_1v2.n31 5.24569
R15662 vbg_1v2.n2 vbg_1v2.n1 4.5005
R15663 vbg_1v2.n4 vbg_1v2.n3 4.5005
R15664 vbg_1v2.n6 vbg_1v2.n5 4.5005
R15665 vbg_1v2.n8 vbg_1v2.n7 4.5005
R15666 vbg_1v2.n10 vbg_1v2.n9 4.5005
R15667 vbg_1v2.n12 vbg_1v2.n11 4.5005
R15668 vbg_1v2.n14 vbg_1v2.n13 4.5005
R15669 vbg_1v2.n16 vbg_1v2.n15 4.5005
R15670 vbg_1v2.n18 vbg_1v2.n17 4.5005
R15671 vbg_1v2.n20 vbg_1v2.n19 4.5005
R15672 vbg_1v2.n22 vbg_1v2.n21 4.5005
R15673 vbg_1v2.n24 vbg_1v2.n23 4.5005
R15674 vbg_1v2.n26 vbg_1v2.n25 4.5005
R15675 vbg_1v2.n28 vbg_1v2.n27 4.5005
R15676 vbg_1v2.n30 vbg_1v2.n29 4.5005
R15677 vbg_1v2.n33 vbg_1v2.n32 4.5005
R15678 vbg_1v2.n35 vbg_1v2.n34 4.5005
R15679 vbg_1v2.n37 vbg_1v2.n36 4.5005
R15680 vbg_1v2.n39 vbg_1v2.n38 4.5005
R15681 vbg_1v2.n41 vbg_1v2.n40 4.5005
R15682 vbg_1v2.n43 vbg_1v2.n42 4.5005
R15683 vbg_1v2.n45 vbg_1v2.n44 4.5005
R15684 vbg_1v2.n47 vbg_1v2.n46 4.5005
R15685 vbg_1v2.n49 vbg_1v2.n48 4.5005
R15686 vbg_1v2.n51 vbg_1v2.n50 4.5005
R15687 vbg_1v2.n53 vbg_1v2.n52 4.5005
R15688 vbg_1v2.n55 vbg_1v2.n54 4.5005
R15689 vbg_1v2.n57 vbg_1v2.n56 4.5005
R15690 vbg_1v2.n59 vbg_1v2.n58 4.5005
R15691 vbg_1v2.n61 vbg_1v2.n60 4.5005
R15692 vbg_1v2.n79 vbg_1v2.n62 4.5005
R15693 vbg_1v2.n81 vbg_1v2.n80 4.5005
R15694 vbg_1v2.n81 vbg_1v2.n62 2.63992
R15695 vbg_1v2.n30 vbg_1v2.n27 0.745692
R15696 vbg_1v2.n26 vbg_1v2.n23 0.745692
R15697 vbg_1v2.n22 vbg_1v2.n19 0.745692
R15698 vbg_1v2.n18 vbg_1v2.n15 0.745692
R15699 vbg_1v2.n14 vbg_1v2.n11 0.745692
R15700 vbg_1v2.n10 vbg_1v2.n7 0.745692
R15701 vbg_1v2.n6 vbg_1v2.n3 0.745692
R15702 vbg_1v2.n61 vbg_1v2.n58 0.745692
R15703 vbg_1v2.n57 vbg_1v2.n54 0.745692
R15704 vbg_1v2.n53 vbg_1v2.n50 0.745692
R15705 vbg_1v2.n49 vbg_1v2.n46 0.745692
R15706 vbg_1v2.n45 vbg_1v2.n42 0.745692
R15707 vbg_1v2.n41 vbg_1v2.n38 0.745692
R15708 vbg_1v2.n37 vbg_1v2.n34 0.745692
R15709 vbg_1v2.n69 vbg_1v2.n68 0.484196
R15710 vbg_1v2.n70 vbg_1v2.n69 0.484196
R15711 vbg_1v2.n70 vbg_1v2.n65 0.484196
R15712 vbg_1v2.n74 vbg_1v2.n65 0.484196
R15713 vbg_1v2.n75 vbg_1v2.n74 0.484196
R15714 vbg_1v2.n76 vbg_1v2.n75 0.484196
R15715 vbg_1v2.n76 vbg_1v2.n63 0.484196
R15716 vbg_1v2.n67 vbg_1v2.n66 0.484196
R15717 vbg_1v2.n71 vbg_1v2.n66 0.484196
R15718 vbg_1v2.n72 vbg_1v2.n71 0.484196
R15719 vbg_1v2.n73 vbg_1v2.n72 0.484196
R15720 vbg_1v2.n73 vbg_1v2.n64 0.484196
R15721 vbg_1v2.n77 vbg_1v2.n64 0.484196
R15722 vbg_1v2.n78 vbg_1v2.n77 0.484196
R15723 vbg_1v2.n80 vbg_1v2.n63 0.459739
R15724 vbg_1v2.n79 vbg_1v2.n78 0.459739
R15725 vbg_1v2.n27 vbg_1v2.n26 0.260115
R15726 vbg_1v2.n23 vbg_1v2.n22 0.260115
R15727 vbg_1v2.n19 vbg_1v2.n18 0.260115
R15728 vbg_1v2.n15 vbg_1v2.n14 0.260115
R15729 vbg_1v2.n11 vbg_1v2.n10 0.260115
R15730 vbg_1v2.n7 vbg_1v2.n6 0.260115
R15731 vbg_1v2.n3 vbg_1v2.n2 0.260115
R15732 vbg_1v2.n58 vbg_1v2.n57 0.260115
R15733 vbg_1v2.n54 vbg_1v2.n53 0.260115
R15734 vbg_1v2.n50 vbg_1v2.n49 0.260115
R15735 vbg_1v2.n46 vbg_1v2.n45 0.260115
R15736 vbg_1v2.n42 vbg_1v2.n41 0.260115
R15737 vbg_1v2.n38 vbg_1v2.n37 0.260115
R15738 vbg_1v2.n34 vbg_1v2.n33 0.260115
R15739 vbg_1v2 vbg_1v2.n81 0.063
R15740 ibias_gen_0.vn0.n9 ibias_gen_0.vn0.t19 50.4613
R15741 ibias_gen_0.vn0.n10 ibias_gen_0.vn0.t19 50.4344
R15742 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.n7 49.6079
R15743 ibias_gen_0.vn0.n4 ibias_gen_0.vn0.t3 49.2687
R15744 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.t3 49.1817
R15745 ibias_gen_0.vn0.t1 ibias_gen_0.vn0.n3 48.1029
R15746 ibias_gen_0.vn0.t20 ibias_gen_0.vn0.n9 48.1029
R15747 ibias_gen_0.vn0.n8 ibias_gen_0.vn0.t1 48.1029
R15748 ibias_gen_0.vn0.n10 ibias_gen_0.vn0.t20 48.1029
R15749 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.t9 22.9447
R15750 ibias_gen_0.Mt4 ibias_gen_0.vn0.n2 21.105
R15751 ibias_gen_0.Mt4 ibias_gen_0.vn0.n15 19.6387
R15752 ibias_gen_0.Mt4 ibias_gen_0.vn0.n14 19.6387
R15753 ibias_gen_0.Mt4 ibias_gen_0.vn0.n13 19.6387
R15754 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.n12 19.6387
R15755 ibias_gen_0.Mt4 ibias_gen_0.vn0.n16 19.6387
R15756 ibias_gen_0.vn0.n6 ibias_gen_0.vn0.n5 13.8791
R15757 ibias_gen_0.vn0.n9 ibias_gen_0.vn0.n8 13.7174
R15758 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.n11 12.7887
R15759 ibias_gen_0.vn0.n11 ibias_gen_0.vn0.n3 7.26784
R15760 ibias_gen_0.vn0.n11 ibias_gen_0.vn0.n10 6.45004
R15761 ibias_gen_0.vn0.n7 ibias_gen_0.vn0.t16 5.5395
R15762 ibias_gen_0.vn0.n7 ibias_gen_0.vn0.t17 5.5395
R15763 ibias_gen_0.vn0.n15 ibias_gen_0.vn0.t8 3.3065
R15764 ibias_gen_0.vn0.n15 ibias_gen_0.vn0.t10 3.3065
R15765 ibias_gen_0.vn0.n14 ibias_gen_0.vn0.t11 3.3065
R15766 ibias_gen_0.vn0.n14 ibias_gen_0.vn0.t13 3.3065
R15767 ibias_gen_0.vn0.n13 ibias_gen_0.vn0.t14 3.3065
R15768 ibias_gen_0.vn0.n13 ibias_gen_0.vn0.t15 3.3065
R15769 ibias_gen_0.vn0.n12 ibias_gen_0.vn0.t6 3.3065
R15770 ibias_gen_0.vn0.n12 ibias_gen_0.vn0.t12 3.3065
R15771 ibias_gen_0.vn0.n5 ibias_gen_0.vn0.t2 3.3065
R15772 ibias_gen_0.vn0.n5 ibias_gen_0.vn0.t4 3.3065
R15773 ibias_gen_0.vn0.n2 ibias_gen_0.vn0.t18 3.3065
R15774 ibias_gen_0.vn0.n2 ibias_gen_0.vn0.t5 3.3065
R15775 ibias_gen_0.vn0.n16 ibias_gen_0.vn0.t0 3.3065
R15776 ibias_gen_0.vn0.n16 ibias_gen_0.vn0.t7 3.3065
R15777 ibias_gen_0.Mt4 ibias_gen_0.vn0.n0 2.11628
R15778 ibias_gen_0.vn0.n6 ibias_gen_0.vn0.n4 1.44615
R15779 ibias_gen_0.vn0.n8 ibias_gen_0.vn0.n1 1.30001
R15780 ibias_gen_0.vn0.n4 ibias_gen_0.vn0.n3 1.16626
R15781 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.n6 1.15267
R15782 ibias_gen_0.vp0.n3 ibias_gen_0.vp0.n1 57.7416
R15783 ibias_gen_0.vp0.n8 ibias_gen_0.vp0.t13 50.9767
R15784 ibias_gen_0.vp0.t13 ibias_gen_0.vp0.n6 50.9767
R15785 ibias_gen_0.vp0.n7 ibias_gen_0.vp0.t8 49.8109
R15786 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.t8 49.7239
R15787 ibias_gen_0.vp0.t10 ibias_gen_0.vp0.n9 48.6451
R15788 ibias_gen_0.vp0.t12 ibias_gen_0.vp0.n6 48.6451
R15789 ibias_gen_0.vp0.n10 ibias_gen_0.vp0.t10 48.6451
R15790 ibias_gen_0.vp0.n8 ibias_gen_0.vp0.t12 48.6451
R15791 ibias_gen_0.vp0.n5 ibias_gen_0.vp0.n4 42.4505
R15792 ibias_gen_0.vp0.n3 ibias_gen_0.vp0.n2 42.4505
R15793 ibias_gen_0.vp0.n14 ibias_gen_0.vp0.n13 18.2113
R15794 ibias_gen_0.vp0.n12 ibias_gen_0.vp0.n11 17.2812
R15795 ibias_gen_0.vp0.n10 ibias_gen_0.vp0.n6 13.7361
R15796 ibias_gen_0.vp0.n9 ibias_gen_0.vp0.n8 13.7361
R15797 ibias_gen_0.vp0.n13 ibias_gen_0.vp0.n12 13.3639
R15798 ibias_gen_0.vp0.n4 ibias_gen_0.vp0.t9 5.5395
R15799 ibias_gen_0.vp0.n4 ibias_gen_0.vp0.t11 5.5395
R15800 ibias_gen_0.vp0.n2 ibias_gen_0.vp0.t7 5.5395
R15801 ibias_gen_0.vp0.n2 ibias_gen_0.vp0.t5 5.5395
R15802 ibias_gen_0.vp0.n1 ibias_gen_0.vp0.t4 5.5395
R15803 ibias_gen_0.vp0.n1 ibias_gen_0.vp0.t6 5.5395
R15804 ibias_gen_0.vp0.n13 ibias_gen_0.vp0.n3 3.97054
R15805 ibias_gen_0.vp0.n12 ibias_gen_0.vp0.n0 3.77198
R15806 ibias_gen_0.vp0.n11 ibias_gen_0.vp0.t2 3.3065
R15807 ibias_gen_0.vp0.n11 ibias_gen_0.vp0.t1 3.3065
R15808 ibias_gen_0.vp0.n14 ibias_gen_0.vp0.t3 3.3065
R15809 ibias_gen_0.vp0.t0 ibias_gen_0.vp0.n14 3.3065
R15810 ibias_gen_0.vp0.n7 ibias_gen_0.vp0.n5 1.47061
R15811 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.n10 1.3293
R15812 ibias_gen_0.vp0.n9 ibias_gen_0.vp0.n7 1.16626
R15813 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.n5 1.13637
R15814 ibias_gen_0.vr.n2 ibias_gen_0.vr.n0 21.7373
R15815 ibias_gen_0.vr.n2 ibias_gen_0.vr.n1 20.4114
R15816 ibias_gen_0.vr.t4 ibias_gen_0.vr.n2 17.6029
R15817 ibias_gen_0.vr.n1 ibias_gen_0.vr.t0 3.3065
R15818 ibias_gen_0.vr.n1 ibias_gen_0.vr.t3 3.3065
R15819 ibias_gen_0.vr.n0 ibias_gen_0.vr.t2 3.3065
R15820 ibias_gen_0.vr.n0 ibias_gen_0.vr.t1 3.3065
R15821 outb.n2 outb.n0 243.458
R15822 outb.n2 outb.n1 205.059
R15823 outb.n4 outb.n3 205.059
R15824 outb.n6 outb.n5 205.059
R15825 outb.n8 outb.n7 205.059
R15826 outb.n10 outb.n9 205.059
R15827 outb.n12 outb.n11 205.059
R15828 outb.n14 outb.n13 205.059
R15829 outb.n17 outb.n15 133.534
R15830 outb.n17 outb.n16 99.1759
R15831 outb.n19 outb.n18 99.1759
R15832 outb.n21 outb.n20 99.1759
R15833 outb.n23 outb.n22 99.1759
R15834 outb.n25 outb.n24 99.1759
R15835 outb.n27 outb.n26 99.1759
R15836 outb outb.n28 97.4305
R15837 outb.n4 outb.n2 38.4005
R15838 outb.n6 outb.n4 38.4005
R15839 outb.n8 outb.n6 38.4005
R15840 outb.n10 outb.n8 38.4005
R15841 outb.n12 outb.n10 38.4005
R15842 outb.n14 outb.n12 38.4005
R15843 outb.n19 outb.n17 34.3584
R15844 outb.n21 outb.n19 34.3584
R15845 outb.n23 outb.n21 34.3584
R15846 outb.n25 outb.n23 34.3584
R15847 outb.n27 outb.n25 34.3584
R15848 outb.n29 outb.n27 34.3584
R15849 outb.n13 outb.t15 26.5955
R15850 outb.n13 outb.t5 26.5955
R15851 outb.n0 outb.t13 26.5955
R15852 outb.n0 outb.t4 26.5955
R15853 outb.n1 outb.t11 26.5955
R15854 outb.n1 outb.t7 26.5955
R15855 outb.n3 outb.t10 26.5955
R15856 outb.n3 outb.t2 26.5955
R15857 outb.n5 outb.t14 26.5955
R15858 outb.n5 outb.t1 26.5955
R15859 outb.n7 outb.t9 26.5955
R15860 outb.n7 outb.t3 26.5955
R15861 outb.n9 outb.t12 26.5955
R15862 outb.n9 outb.t8 26.5955
R15863 outb.n11 outb.t0 26.5955
R15864 outb.n11 outb.t6 26.5955
R15865 outb.n28 outb.t28 24.9236
R15866 outb.n28 outb.t18 24.9236
R15867 outb.n15 outb.t26 24.9236
R15868 outb.n15 outb.t17 24.9236
R15869 outb.n16 outb.t24 24.9236
R15870 outb.n16 outb.t20 24.9236
R15871 outb.n18 outb.t23 24.9236
R15872 outb.n18 outb.t31 24.9236
R15873 outb.n20 outb.t27 24.9236
R15874 outb.n20 outb.t30 24.9236
R15875 outb.n22 outb.t22 24.9236
R15876 outb.n22 outb.t16 24.9236
R15877 outb.n24 outb.t25 24.9236
R15878 outb.n24 outb.t21 24.9236
R15879 outb.n26 outb.t29 24.9236
R15880 outb.n26 outb.t19 24.9236
R15881 outb outb.n14 18.4247
R15882 outb.n30 outb.n29 10.0853
R15883 outb.n30 outb 4.84706
R15884 outb.n29 outb 1.74595
R15885 outb outb.n30 1.35808
R15886 ibias_gen_0.vp.n10 ibias_gen_0.vp.t4 56.5501
R15887 ibias_gen_0.vp.n4 ibias_gen_0.vp.t11 50.9767
R15888 ibias_gen_0.vp.n5 ibias_gen_0.vp.t11 50.9767
R15889 ibias_gen_0.vp.t9 ibias_gen_0.vp.n6 50.9767
R15890 ibias_gen_0.vp.t8 ibias_gen_0.vp.n4 48.6451
R15891 ibias_gen_0.vp.n7 ibias_gen_0.vp.t9 48.6451
R15892 ibias_gen_0.vp.n6 ibias_gen_0.vp.t7 48.6451
R15893 ibias_gen_0.vp.n5 ibias_gen_0.vp.t8 48.6451
R15894 ibias_gen_0.vp.t7 ibias_gen_0.vp.n3 48.6451
R15895 ibias_gen_0.vp.n0 ibias_gen_0.vp.n11 42.5266
R15896 ibias_gen_0.vp.n0 ibias_gen_0.vp.n2 42.4505
R15897 ibias_gen_0.vp.n9 ibias_gen_0.vp.n8 26.1532
R15898 ibias_gen_0.vp.n8 ibias_gen_0.vp.t12 25.4891
R15899 ibias_gen_0.vp.n8 ibias_gen_0.vp.t10 24.3233
R15900 ibias_gen_0.vp.n13 ibias_gen_0.vp.n12 15.1165
R15901 ibias_gen_0.vp.n12 ibias_gen_0.vp.n1 14.8365
R15902 ibias_gen_0.vp.n10 ibias_gen_0.vp.n9 8.08875
R15903 ibias_gen_0.vp.n12 ibias_gen_0.vp.n0 7.57893
R15904 ibias_gen_0.vp.n0 ibias_gen_0.vp.n10 6.28836
R15905 ibias_gen_0.vp.n2 ibias_gen_0.vp.t1 5.5395
R15906 ibias_gen_0.vp.t3 ibias_gen_0.vp.n2 5.5395
R15907 ibias_gen_0.vp.n11 ibias_gen_0.vp.t3 5.5395
R15908 ibias_gen_0.vp.n11 ibias_gen_0.vp.t6 5.5395
R15909 ibias_gen_0.vp.n1 ibias_gen_0.vp.t5 3.3065
R15910 ibias_gen_0.vp.t0 ibias_gen_0.vp.n1 3.3065
R15911 ibias_gen_0.vp.t0 ibias_gen_0.vp.n13 3.3065
R15912 ibias_gen_0.vp.n13 ibias_gen_0.vp.t2 3.3065
R15913 ibias_gen_0.vp.n9 ibias_gen_0.vp.n7 2.37524
R15914 ibias_gen_0.vp.n6 ibias_gen_0.vp.n5 2.33202
R15915 ibias_gen_0.vp.n4 ibias_gen_0.vp.n3 2.33202
R15916 ibias_gen_0.vp.n7 ibias_gen_0.vp.n3 2.33126
R15917 itest itest.n0 45.907
R15918 itest.n0 itest.t0 5.5395
R15919 itest.n0 itest.t1 5.5395
R15920 rstring_mux_0.vtrip7.n5 rstring_mux_0.vtrip7.n3 50.7022
R15921 rstring_mux_0.vtrip7.n2 rstring_mux_0.vtrip7.n0 50.7022
R15922 rstring_mux_0.vtrip7.n6 rstring_mux_0.vtrip7.n5 15.3935
R15923 rstring_mux_0.vtrip7.n5 rstring_mux_0.vtrip7.n4 13.8791
R15924 rstring_mux_0.vtrip7.n2 rstring_mux_0.vtrip7.n1 13.8791
R15925 rstring_mux_0.vtrip7.t0 rstring_mux_0.vtrip7.n7 10.5857
R15926 rstring_mux_0.vtrip7.n7 rstring_mux_0.vtrip7.t1 10.5847
R15927 rstring_mux_0.vtrip7.n3 rstring_mux_0.vtrip7.t5 5.5395
R15928 rstring_mux_0.vtrip7.n3 rstring_mux_0.vtrip7.t4 5.5395
R15929 rstring_mux_0.vtrip7.n0 rstring_mux_0.vtrip7.t2 5.5395
R15930 rstring_mux_0.vtrip7.n0 rstring_mux_0.vtrip7.t3 5.5395
R15931 rstring_mux_0.vtrip7.n6 rstring_mux_0.vtrip7.n2 5.2741
R15932 rstring_mux_0.vtrip7.n4 rstring_mux_0.vtrip7.t6 3.3065
R15933 rstring_mux_0.vtrip7.n4 rstring_mux_0.vtrip7.t7 3.3065
R15934 rstring_mux_0.vtrip7.n1 rstring_mux_0.vtrip7.t8 3.3065
R15935 rstring_mux_0.vtrip7.n1 rstring_mux_0.vtrip7.t9 3.3065
R15936 rstring_mux_0.vtrip7.n7 rstring_mux_0.vtrip7.n6 2.48711
R15937 rstring_mux_0.vtrip2.n5 rstring_mux_0.vtrip2.n3 50.7022
R15938 rstring_mux_0.vtrip2.n2 rstring_mux_0.vtrip2.n0 50.7022
R15939 rstring_mux_0.vtrip2.n7 rstring_mux_0.vtrip2.n6 23.8383
R15940 rstring_mux_0.vtrip2.n6 rstring_mux_0.vtrip2.n5 14.3726
R15941 rstring_mux_0.vtrip2.n5 rstring_mux_0.vtrip2.n4 13.8791
R15942 rstring_mux_0.vtrip2.n2 rstring_mux_0.vtrip2.n1 13.8791
R15943 rstring_mux_0.vtrip2.n7 rstring_mux_0.vtrip2.t3 10.6303
R15944 rstring_mux_0.vtrip2.n3 rstring_mux_0.vtrip2.t7 5.5395
R15945 rstring_mux_0.vtrip2.n3 rstring_mux_0.vtrip2.t6 5.5395
R15946 rstring_mux_0.vtrip2.n0 rstring_mux_0.vtrip2.t0 5.5395
R15947 rstring_mux_0.vtrip2.n0 rstring_mux_0.vtrip2.t1 5.5395
R15948 rstring_mux_0.vtrip2.n6 rstring_mux_0.vtrip2.n2 4.21994
R15949 rstring_mux_0.vtrip2.n4 rstring_mux_0.vtrip2.t8 3.3065
R15950 rstring_mux_0.vtrip2.n4 rstring_mux_0.vtrip2.t9 3.3065
R15951 rstring_mux_0.vtrip2.n1 rstring_mux_0.vtrip2.t5 3.3065
R15952 rstring_mux_0.vtrip2.n1 rstring_mux_0.vtrip2.t4 3.3065
R15953 rstring_mux_0.vtrip2 rstring_mux_0.vtrip2.t2 0.769662
R15954 rstring_mux_0.vtrip2 rstring_mux_0.vtrip2.n7 0.0563195
R15955 ibias_gen_0.vp1.n5 ibias_gen_0.vp1.n4 53.0003
R15956 ibias_gen_0.vp1.t8 ibias_gen_0.vp1.n3 49.8109
R15957 ibias_gen_0.vp1.n3 ibias_gen_0.vp1.t6 49.8109
R15958 ibias_gen_0.vp1.t6 ibias_gen_0.vp1.n0 49.7878
R15959 ibias_gen_0.vp1.n0 ibias_gen_0.vp1.t8 49.6053
R15960 ibias_gen_0.vp1 ibias_gen_0.vp1.n6 45.7548
R15961 ibias_gen_0.vp1.n2 ibias_gen_0.vp1.n1 42.4505
R15962 ibias_gen_0.vp1.n9 ibias_gen_0.vp1.n7 18.5825
R15963 ibias_gen_0.vp1.n15 ibias_gen_0.vp1.n14 17.1535
R15964 ibias_gen_0.vp1.n11 ibias_gen_0.vp1.n10 16.3247
R15965 ibias_gen_0.vp1.n9 ibias_gen_0.vp1.n8 16.3247
R15966 ibias_gen_0.vp1.n13 ibias_gen_0.vp1.n12 15.5548
R15967 ibias_gen_0.vp1.n15 ibias_gen_0.vp1.n13 11.684
R15968 ibias_gen_0.vp1.n6 ibias_gen_0.vp1.t11 5.5395
R15969 ibias_gen_0.vp1.n6 ibias_gen_0.vp1.t10 5.5395
R15970 ibias_gen_0.vp1.n4 ibias_gen_0.vp1.t15 5.5395
R15971 ibias_gen_0.vp1.n4 ibias_gen_0.vp1.t17 5.5395
R15972 ibias_gen_0.vp1.n1 ibias_gen_0.vp1.t7 5.5395
R15973 ibias_gen_0.vp1.n1 ibias_gen_0.vp1.t9 5.5395
R15974 ibias_gen_0.vp1.n5 ibias_gen_0.vp1.n0 4.85318
R15975 ibias_gen_0.vp1.n11 ibias_gen_0.vp1.n9 4.51612
R15976 ibias_gen_0.vp1.n12 ibias_gen_0.vp1.t12 3.3065
R15977 ibias_gen_0.vp1.n12 ibias_gen_0.vp1.t1 3.3065
R15978 ibias_gen_0.vp1.n10 ibias_gen_0.vp1.t14 3.3065
R15979 ibias_gen_0.vp1.n10 ibias_gen_0.vp1.t5 3.3065
R15980 ibias_gen_0.vp1.n8 ibias_gen_0.vp1.t4 3.3065
R15981 ibias_gen_0.vp1.n8 ibias_gen_0.vp1.t13 3.3065
R15982 ibias_gen_0.vp1.n7 ibias_gen_0.vp1.t2 3.3065
R15983 ibias_gen_0.vp1.n7 ibias_gen_0.vp1.t3 3.3065
R15984 ibias_gen_0.vp1.n14 ibias_gen_0.vp1.t0 3.3065
R15985 ibias_gen_0.vp1.n14 ibias_gen_0.vp1.t16 3.3065
R15986 ibias_gen_0.vp1.n13 ibias_gen_0.vp1.n11 2.27562
R15987 ibias_gen_0.vp1 ibias_gen_0.vp1.n15 1.87819
R15988 ibias_gen_0.vp1.n2 ibias_gen_0.vp1.n0 1.48628
R15989 ibias_gen_0.vp1.n3 ibias_gen_0.vp1.n2 1.47061
R15990 ibias_gen_0.vp1 ibias_gen_0.vp1.n5 1.36236
R15991 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n1 47.4959
R15992 ibias_gen_0.vn1.n3 ibias_gen_0.vn1.t14 27.5855
R15993 ibias_gen_0.vn1.n2 ibias_gen_0.vn1.t10 27.5855
R15994 ibias_gen_0.vn1.n6 ibias_gen_0.vn1.t16 27.5855
R15995 ibias_gen_0.vn1.n5 ibias_gen_0.vn1.t12 27.5855
R15996 ibias_gen_0.vn1.n10 ibias_gen_0.vn1.t3 26.004
R15997 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n13 24.5059
R15998 ibias_gen_0.vn1.n3 ibias_gen_0.vn1.t17 24.3247
R15999 ibias_gen_0.vn1.n2 ibias_gen_0.vn1.t15 24.3247
R16000 ibias_gen_0.vn1.n6 ibias_gen_0.vn1.t13 24.3247
R16001 ibias_gen_0.vn1.n5 ibias_gen_0.vn1.t11 24.3247
R16002 ibias_gen_0.vn1.n9 ibias_gen_0.vn1.t1 24.3247
R16003 ibias_gen_0.vn1.n14 ibias_gen_0.vn1.n0 17.1535
R16004 ibias_gen_0.vn1.n12 ibias_gen_0.vn1.n11 13.8791
R16005 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n12 12.7397
R16006 ibias_gen_0.vn1.n1 ibias_gen_0.vn1.t7 5.5395
R16007 ibias_gen_0.vn1.n1 ibias_gen_0.vn1.t8 5.5395
R16008 ibias_gen_0.vn1.n4 ibias_gen_0.vn1.n2 4.66645
R16009 ibias_gen_0.vn1.n7 ibias_gen_0.vn1.n5 4.66645
R16010 ibias_gen_0.vn1.n13 ibias_gen_0.vn1.t5 3.3065
R16011 ibias_gen_0.vn1.n13 ibias_gen_0.vn1.t6 3.3065
R16012 ibias_gen_0.vn1.n11 ibias_gen_0.vn1.t2 3.3065
R16013 ibias_gen_0.vn1.n11 ibias_gen_0.vn1.t4 3.3065
R16014 ibias_gen_0.vn1.n14 ibias_gen_0.vn1.t9 3.3065
R16015 ibias_gen_0.vn1.t0 ibias_gen_0.vn1.n14 3.3065
R16016 ibias_gen_0.vn1.n8 ibias_gen_0.vn1.n4 2.41645
R16017 ibias_gen_0.vn1.n8 ibias_gen_0.vn1.n7 2.41645
R16018 ibias_gen_0.vn1.n4 ibias_gen_0.vn1.n3 2.2505
R16019 ibias_gen_0.vn1.n7 ibias_gen_0.vn1.n6 2.2505
R16020 ibias_gen_0.vn1.n9 ibias_gen_0.vn1.n8 2.2505
R16021 ibias_gen_0.vn1.n10 ibias_gen_0.vn1.n9 1.58202
R16022 ibias_gen_0.vn1.n12 ibias_gen_0.vn1.n10 1.37822
R16023 vtrip_decoded[3].n0 vtrip_decoded[3].t1 186.374
R16024 vtrip_decoded[3].n0 vtrip_decoded[3].t0 170.308
R16025 vtrip_decoded[3] vtrip_decoded[3].n1 154.56
R16026 vtrip_decoded[3].n2 vtrip_decoded[3].n1 153.462
R16027 vtrip_decoded[3].n1 vtrip_decoded[3].n0 101.513
R16028 vtrip_decoded[3].n3 vtrip_decoded[3] 11.8005
R16029 vtrip_decoded[3].n3 vtrip_decoded[3].n2 4.96991
R16030 vtrip_decoded[3].n2 vtrip_decoded[3] 3.46403
R16031 vtrip_decoded[3] vtrip_decoded[3].n3 2.71109
R16032 osc_ena.n1 osc_ena.t3 413.582
R16033 osc_ena.n0 osc_ena.t0 348.789
R16034 osc_ena.n1 osc_ena.t1 227.718
R16035 osc_ena.n0 osc_ena.t2 224.327
R16036 osc_ena.n2 osc_ena.n0 13.8663
R16037 osc_ena.n2 osc_ena.n1 4.5005
R16038 osc_ena osc_ena.n2 0.0755
R16039 rstring_mux_0.vtrip3.n5 rstring_mux_0.vtrip3.n3 50.7022
R16040 rstring_mux_0.vtrip3.n2 rstring_mux_0.vtrip3.n0 50.7022
R16041 rstring_mux_0.vtrip3.n6 rstring_mux_0.vtrip3.n5 14.2209
R16042 rstring_mux_0.vtrip3.n5 rstring_mux_0.vtrip3.n4 13.8791
R16043 rstring_mux_0.vtrip3.n2 rstring_mux_0.vtrip3.n1 13.8791
R16044 rstring_mux_0.vtrip3.t0 rstring_mux_0.vtrip3.n7 10.5857
R16045 rstring_mux_0.vtrip3.n7 rstring_mux_0.vtrip3.t9 10.5847
R16046 rstring_mux_0.vtrip3.n6 rstring_mux_0.vtrip3.n2 5.7125
R16047 rstring_mux_0.vtrip3.n3 rstring_mux_0.vtrip3.t5 5.5395
R16048 rstring_mux_0.vtrip3.n3 rstring_mux_0.vtrip3.t6 5.5395
R16049 rstring_mux_0.vtrip3.n0 rstring_mux_0.vtrip3.t3 5.5395
R16050 rstring_mux_0.vtrip3.n0 rstring_mux_0.vtrip3.t4 5.5395
R16051 rstring_mux_0.vtrip3.n4 rstring_mux_0.vtrip3.t2 3.3065
R16052 rstring_mux_0.vtrip3.n4 rstring_mux_0.vtrip3.t1 3.3065
R16053 rstring_mux_0.vtrip3.n1 rstring_mux_0.vtrip3.t7 3.3065
R16054 rstring_mux_0.vtrip3.n1 rstring_mux_0.vtrip3.t8 3.3065
R16055 rstring_mux_0.vtrip3.n7 rstring_mux_0.vtrip3.n6 3.16869
R16056 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.t0 56.685
R16057 ibias_gen_0.vstart.n5 ibias_gen_0.vstart.n3 20.328
R16058 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.n1 20.2356
R16059 ibias_gen_0.vstart.n5 ibias_gen_0.vstart.n4 20.069
R16060 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.n2 20.069
R16061 ibias_gen_0.vstart.n7 ibias_gen_0.vstart.n6 20.069
R16062 ibias_gen_0.vstart.n4 ibias_gen_0.vstart.t10 3.3065
R16063 ibias_gen_0.vstart.n4 ibias_gen_0.vstart.t1 3.3065
R16064 ibias_gen_0.vstart.n3 ibias_gen_0.vstart.t7 3.3065
R16065 ibias_gen_0.vstart.n3 ibias_gen_0.vstart.t4 3.3065
R16066 ibias_gen_0.vstart.n2 ibias_gen_0.vstart.t5 3.3065
R16067 ibias_gen_0.vstart.n2 ibias_gen_0.vstart.t6 3.3065
R16068 ibias_gen_0.vstart.n1 ibias_gen_0.vstart.t2 3.3065
R16069 ibias_gen_0.vstart.n1 ibias_gen_0.vstart.t3 3.3065
R16070 ibias_gen_0.vstart.n7 ibias_gen_0.vstart.t8 3.3065
R16071 ibias_gen_0.vstart.t9 ibias_gen_0.vstart.n7 3.3065
R16072 ibias_gen_0.vstart.n6 ibias_gen_0.vstart.n0 0.280933
R16073 ibias_gen_0.vstart.n6 ibias_gen_0.vstart.n5 0.2449
R16074 schmitt_trigger_0.out.n8 schmitt_trigger_0.out.t12 248.236
R16075 schmitt_trigger_0.out.n6 schmitt_trigger_0.out.t11 240.778
R16076 schmitt_trigger_0.out.n7 schmitt_trigger_0.out.t4 240.613
R16077 schmitt_trigger_0.out.n6 schmitt_trigger_0.out.t5 240.349
R16078 schmitt_trigger_0.out.n5 schmitt_trigger_0.out.t1 236.369
R16079 schmitt_trigger_0.out.n0 schmitt_trigger_0.out.t8 212.081
R16080 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.t7 212.081
R16081 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.t13 212.081
R16082 schmitt_trigger_0.out.n3 schmitt_trigger_0.out.t6 212.081
R16083 schmitt_trigger_0.out.n5 schmitt_trigger_0.out.n4 207.585
R16084 schmitt_trigger_0.out.n12 schmitt_trigger_0.out.n3 188.516
R16085 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n1 154.304
R16086 schmitt_trigger_0.out.n14 schmitt_trigger_0.out.n13 152
R16087 schmitt_trigger_0.out.n17 schmitt_trigger_0.out.n16 152
R16088 schmitt_trigger_0.out.n0 schmitt_trigger_0.out.t14 139.78
R16089 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.t10 139.78
R16090 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.t15 139.78
R16091 schmitt_trigger_0.out.n3 schmitt_trigger_0.out.t9 139.78
R16092 schmitt_trigger_0.out.n10 schmitt_trigger_0.out.t3 91.727
R16093 schmitt_trigger_0.out.n1 schmitt_trigger_0.out.n0 30.6732
R16094 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.n1 30.6732
R16095 schmitt_trigger_0.out.n16 schmitt_trigger_0.out.n2 30.6732
R16096 schmitt_trigger_0.out.n16 schmitt_trigger_0.out.n15 30.6732
R16097 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.n14 30.6732
R16098 schmitt_trigger_0.out.n14 schmitt_trigger_0.out.n3 30.6732
R16099 schmitt_trigger_0.out.n4 schmitt_trigger_0.out.t2 28.5655
R16100 schmitt_trigger_0.out.n4 schmitt_trigger_0.out.t0 28.5655
R16101 schmitt_trigger_0.out.n11 schmitt_trigger_0.out.n10 20.1312
R16102 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n17 19.2005
R16103 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n12 17.1525
R16104 schmitt_trigger_0.out.n11 sky130_fd_sc_hd__inv_4_0.A 12.8005
R16105 schmitt_trigger_0.out.n9 schmitt_trigger_0.out.n5 8.66251
R16106 schmitt_trigger_0.out.n13 sky130_fd_sc_hd__inv_4_0.A 6.4005
R16107 schmitt_trigger_0.out.n12 sky130_fd_sc_hd__inv_4_0.A 6.4005
R16108 schmitt_trigger_0.out.n8 schmitt_trigger_0.out.n7 4.94425
R16109 schmitt_trigger_0.out.n17 sky130_fd_sc_hd__inv_4_0.A 4.3525
R16110 schmitt_trigger_0.out.n13 schmitt_trigger_0.out.n11 4.3525
R16111 schmitt_trigger_0.out.n9 schmitt_trigger_0.out.n8 4.05633
R16112 schmitt_trigger_0.out.n10 schmitt_trigger_0.out.n9 0.230017
R16113 schmitt_trigger_0.out.n7 schmitt_trigger_0.out.n6 0.117348
R16114 otrip_decoded[6].n0 otrip_decoded[6].t0 186.374
R16115 otrip_decoded[6].n0 otrip_decoded[6].t1 170.308
R16116 otrip_decoded[6] otrip_decoded[6].n1 154.56
R16117 otrip_decoded[6].n2 otrip_decoded[6].n1 153.462
R16118 otrip_decoded[6].n1 otrip_decoded[6].n0 101.513
R16119 otrip_decoded[6].n3 otrip_decoded[6] 11.8005
R16120 otrip_decoded[6].n3 otrip_decoded[6].n2 4.96991
R16121 otrip_decoded[6].n2 otrip_decoded[6] 3.46403
R16122 otrip_decoded[6] otrip_decoded[6].n3 2.71109
R16123 rstring_mux_0.vtrip5.n5 rstring_mux_0.vtrip5.n3 50.7022
R16124 rstring_mux_0.vtrip5.n2 rstring_mux_0.vtrip5.n0 50.7022
R16125 rstring_mux_0.vtrip5.n6 rstring_mux_0.vtrip5.n2 14.7069
R16126 rstring_mux_0.vtrip5.n5 rstring_mux_0.vtrip5.n4 13.8791
R16127 rstring_mux_0.vtrip5.n2 rstring_mux_0.vtrip5.n1 13.8791
R16128 rstring_mux_0.vtrip5.t8 rstring_mux_0.vtrip5.n7 10.5857
R16129 rstring_mux_0.vtrip5.n7 rstring_mux_0.vtrip5.t9 10.5847
R16130 rstring_mux_0.vtrip5.n3 rstring_mux_0.vtrip5.t4 5.5395
R16131 rstring_mux_0.vtrip5.n3 rstring_mux_0.vtrip5.t5 5.5395
R16132 rstring_mux_0.vtrip5.n0 rstring_mux_0.vtrip5.t7 5.5395
R16133 rstring_mux_0.vtrip5.n0 rstring_mux_0.vtrip5.t6 5.5395
R16134 rstring_mux_0.vtrip5.n7 rstring_mux_0.vtrip5.n6 5.07153
R16135 rstring_mux_0.vtrip5.n6 rstring_mux_0.vtrip5.n5 3.33746
R16136 rstring_mux_0.vtrip5.n4 rstring_mux_0.vtrip5.t2 3.3065
R16137 rstring_mux_0.vtrip5.n4 rstring_mux_0.vtrip5.t3 3.3065
R16138 rstring_mux_0.vtrip5.n1 rstring_mux_0.vtrip5.t1 3.3065
R16139 rstring_mux_0.vtrip5.n1 rstring_mux_0.vtrip5.t0 3.3065
R16140 outb_unbuf.n2 outb_unbuf.t3 212.081
R16141 outb_unbuf.n1 outb_unbuf.t2 212.081
R16142 outb_unbuf.n6 outb_unbuf.t6 212.081
R16143 outb_unbuf.n8 outb_unbuf.t1 212.081
R16144 outb_unbuf.n9 outb_unbuf.n8 188.516
R16145 outb_unbuf outb_unbuf.n3 154.304
R16146 outb_unbuf.n5 outb_unbuf.n4 152
R16147 outb_unbuf.n7 outb_unbuf.n0 152
R16148 outb_unbuf.n2 outb_unbuf.t7 139.78
R16149 outb_unbuf.n1 outb_unbuf.t5 139.78
R16150 outb_unbuf.n6 outb_unbuf.t0 139.78
R16151 outb_unbuf.n8 outb_unbuf.t4 139.78
R16152 outb_unbuf.n3 outb_unbuf.n2 30.6732
R16153 outb_unbuf.n3 outb_unbuf.n1 30.6732
R16154 outb_unbuf.n5 outb_unbuf.n1 30.6732
R16155 outb_unbuf.n6 outb_unbuf.n5 30.6732
R16156 outb_unbuf.n7 outb_unbuf.n6 30.6732
R16157 outb_unbuf.n8 outb_unbuf.n7 30.6732
R16158 outb_unbuf.n4 outb_unbuf 19.2005
R16159 outb_unbuf.n10 outb_unbuf 17.3413
R16160 outb_unbuf outb_unbuf.n0 17.1525
R16161 outb_unbuf outb_unbuf.n10 12.5445
R16162 outb_unbuf outb_unbuf.n0 6.4005
R16163 outb_unbuf.n9 outb_unbuf 6.4005
R16164 outb_unbuf.n10 outb_unbuf.n9 4.6085
R16165 outb_unbuf.n4 outb_unbuf 4.3525
R16166 otrip_decoded[4].n0 otrip_decoded[4].t0 186.374
R16167 otrip_decoded[4].n0 otrip_decoded[4].t1 170.308
R16168 otrip_decoded[4] otrip_decoded[4].n1 154.56
R16169 otrip_decoded[4].n2 otrip_decoded[4].n1 153.462
R16170 otrip_decoded[4].n1 otrip_decoded[4].n0 101.513
R16171 otrip_decoded[4].n3 otrip_decoded[4] 11.8005
R16172 otrip_decoded[4].n3 otrip_decoded[4].n2 4.96991
R16173 otrip_decoded[4].n2 otrip_decoded[4] 3.46403
R16174 otrip_decoded[4] otrip_decoded[4].n3 2.71109
R16175 vtrip_decoded[1].n0 vtrip_decoded[1].t1 186.374
R16176 vtrip_decoded[1].n0 vtrip_decoded[1].t0 170.308
R16177 vtrip_decoded[1] vtrip_decoded[1].n1 154.56
R16178 vtrip_decoded[1].n2 vtrip_decoded[1].n1 153.462
R16179 vtrip_decoded[1].n1 vtrip_decoded[1].n0 101.513
R16180 vtrip_decoded[1].n3 vtrip_decoded[1] 11.8005
R16181 vtrip_decoded[1].n3 vtrip_decoded[1].n2 4.96991
R16182 vtrip_decoded[1].n2 vtrip_decoded[1] 3.46403
R16183 vtrip_decoded[1] vtrip_decoded[1].n3 2.71109
R16184 rstring_mux_0.vtrip1.n5 rstring_mux_0.vtrip1.n3 50.7022
R16185 rstring_mux_0.vtrip1.n2 rstring_mux_0.vtrip1.n0 50.7022
R16186 rstring_mux_0.vtrip1.n6 rstring_mux_0.vtrip1.n5 14.0767
R16187 rstring_mux_0.vtrip1.n5 rstring_mux_0.vtrip1.n4 13.8791
R16188 rstring_mux_0.vtrip1.n2 rstring_mux_0.vtrip1.n1 13.8791
R16189 rstring_mux_0.vtrip1.t0 rstring_mux_0.vtrip1.n7 10.5857
R16190 rstring_mux_0.vtrip1.n7 rstring_mux_0.vtrip1.t7 10.5847
R16191 rstring_mux_0.vtrip1.n7 rstring_mux_0.vtrip1.n6 5.61984
R16192 rstring_mux_0.vtrip1.n3 rstring_mux_0.vtrip1.t2 5.5395
R16193 rstring_mux_0.vtrip1.n3 rstring_mux_0.vtrip1.t1 5.5395
R16194 rstring_mux_0.vtrip1.n0 rstring_mux_0.vtrip1.t6 5.5395
R16195 rstring_mux_0.vtrip1.n0 rstring_mux_0.vtrip1.t5 5.5395
R16196 rstring_mux_0.vtrip1.n6 rstring_mux_0.vtrip1.n2 3.9186
R16197 rstring_mux_0.vtrip1.n4 rstring_mux_0.vtrip1.t8 3.3065
R16198 rstring_mux_0.vtrip1.n4 rstring_mux_0.vtrip1.t9 3.3065
R16199 rstring_mux_0.vtrip1.n1 rstring_mux_0.vtrip1.t4 3.3065
R16200 rstring_mux_0.vtrip1.n1 rstring_mux_0.vtrip1.t3 3.3065
R16201 otrip_decoded[2].n0 otrip_decoded[2].t0 186.374
R16202 otrip_decoded[2].n0 otrip_decoded[2].t1 170.308
R16203 otrip_decoded[2] otrip_decoded[2].n1 154.56
R16204 otrip_decoded[2].n2 otrip_decoded[2].n1 153.462
R16205 otrip_decoded[2].n1 otrip_decoded[2].n0 101.513
R16206 otrip_decoded[2].n3 otrip_decoded[2] 11.8005
R16207 otrip_decoded[2].n3 otrip_decoded[2].n2 4.96991
R16208 otrip_decoded[2].n2 otrip_decoded[2] 3.46403
R16209 otrip_decoded[2] otrip_decoded[2].n3 2.71109
R16210 rstring_mux_0.vtrip6.n5 rstring_mux_0.vtrip6.n3 50.7022
R16211 rstring_mux_0.vtrip6.n2 rstring_mux_0.vtrip6.n0 50.7022
R16212 rstring_mux_0.vtrip6.n7 rstring_mux_0.vtrip6.n6 21.6754
R16213 rstring_mux_0.vtrip6.n6 rstring_mux_0.vtrip6.n5 14.944
R16214 rstring_mux_0.vtrip6.n5 rstring_mux_0.vtrip6.n4 13.8791
R16215 rstring_mux_0.vtrip6.n2 rstring_mux_0.vtrip6.n1 13.8791
R16216 rstring_mux_0.vtrip6.n7 rstring_mux_0.vtrip6.t5 10.6303
R16217 rstring_mux_0.vtrip6.n3 rstring_mux_0.vtrip6.t2 5.5395
R16218 rstring_mux_0.vtrip6.n3 rstring_mux_0.vtrip6.t1 5.5395
R16219 rstring_mux_0.vtrip6.n0 rstring_mux_0.vtrip6.t7 5.5395
R16220 rstring_mux_0.vtrip6.n0 rstring_mux_0.vtrip6.t6 5.5395
R16221 rstring_mux_0.vtrip6.n6 rstring_mux_0.vtrip6.n2 5.01904
R16222 rstring_mux_0.vtrip6.n4 rstring_mux_0.vtrip6.t9 3.3065
R16223 rstring_mux_0.vtrip6.n4 rstring_mux_0.vtrip6.t8 3.3065
R16224 rstring_mux_0.vtrip6.n1 rstring_mux_0.vtrip6.t4 3.3065
R16225 rstring_mux_0.vtrip6.n1 rstring_mux_0.vtrip6.t3 3.3065
R16226 rstring_mux_0.vtrip6 rstring_mux_0.vtrip6.t0 0.769662
R16227 rstring_mux_0.vtrip6 rstring_mux_0.vtrip6.n7 0.0563195
R16228 ibias_gen_0.ve.t1 ibias_gen_0.ve.n0 31121.7
R16229 ibias_gen_0.ve.n1 ibias_gen_0.ve.t1 146.25
R16230 ibias_gen_0.ve.n5 ibias_gen_0.ve.n4 62.2607
R16231 ibias_gen_0.ve.n4 ibias_gen_0.ve.n3 21.4545
R16232 ibias_gen_0.ve.n4 ibias_gen_0.ve.n2 20.7025
R16233 ibias_gen_0.ve.n5 ibias_gen_0.ve.n1 8.57525
R16234 sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter ibias_gen_0.ve.n5 6.71196
R16235 ibias_gen_0.ve.n3 ibias_gen_0.ve.t4 3.3065
R16236 ibias_gen_0.ve.n3 ibias_gen_0.ve.t0 3.3065
R16237 ibias_gen_0.ve.n2 ibias_gen_0.ve.t2 3.3065
R16238 ibias_gen_0.ve.n2 ibias_gen_0.ve.t3 3.3065
R16239 sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter ibias_gen_0.ve.n1 1.86379
R16240 rstring_mux_0.vtrip0.n5 rstring_mux_0.vtrip0.n3 50.7022
R16241 rstring_mux_0.vtrip0.n2 rstring_mux_0.vtrip0.n0 50.7022
R16242 rstring_mux_0.vtrip0.n7 rstring_mux_0.vtrip0.n6 25.1771
R16243 rstring_mux_0.vtrip0.n5 rstring_mux_0.vtrip0.n4 13.8791
R16244 rstring_mux_0.vtrip0.n2 rstring_mux_0.vtrip0.n1 13.8791
R16245 rstring_mux_0.vtrip0.n6 rstring_mux_0.vtrip0.n5 13.7519
R16246 rstring_mux_0.vtrip0 rstring_mux_0.vtrip0.t5 10.5739
R16247 rstring_mux_0.vtrip0.n3 rstring_mux_0.vtrip0.t4 5.5395
R16248 rstring_mux_0.vtrip0.n3 rstring_mux_0.vtrip0.t3 5.5395
R16249 rstring_mux_0.vtrip0.n0 rstring_mux_0.vtrip0.t1 5.5395
R16250 rstring_mux_0.vtrip0.n0 rstring_mux_0.vtrip0.t2 5.5395
R16251 rstring_mux_0.vtrip0.n6 rstring_mux_0.vtrip0.n2 3.60196
R16252 rstring_mux_0.vtrip0.n4 rstring_mux_0.vtrip0.t8 3.3065
R16253 rstring_mux_0.vtrip0.n4 rstring_mux_0.vtrip0.t9 3.3065
R16254 rstring_mux_0.vtrip0.n1 rstring_mux_0.vtrip0.t7 3.3065
R16255 rstring_mux_0.vtrip0.n1 rstring_mux_0.vtrip0.t6 3.3065
R16256 rstring_mux_0.vtrip0.n7 rstring_mux_0.vtrip0.t0 0.826075
R16257 rstring_mux_0.vtrip0 rstring_mux_0.vtrip0.n7 0.0563195
R16258 vtrip_decoded[2].n0 vtrip_decoded[2].t1 186.374
R16259 vtrip_decoded[2].n0 vtrip_decoded[2].t0 170.308
R16260 vtrip_decoded[2] vtrip_decoded[2].n1 154.56
R16261 vtrip_decoded[2].n2 vtrip_decoded[2].n1 153.462
R16262 vtrip_decoded[2].n1 vtrip_decoded[2].n0 101.513
R16263 vtrip_decoded[2].n3 vtrip_decoded[2] 11.8005
R16264 vtrip_decoded[2].n3 vtrip_decoded[2].n2 4.96991
R16265 vtrip_decoded[2].n2 vtrip_decoded[2] 3.46403
R16266 vtrip_decoded[2] vtrip_decoded[2].n3 2.71109
R16267 isrc_sel.n0 isrc_sel.t1 186.374
R16268 isrc_sel.n0 isrc_sel.t0 170.308
R16269 isrc_sel isrc_sel.n1 154.56
R16270 isrc_sel.n2 isrc_sel.n1 153.462
R16271 isrc_sel.n1 isrc_sel.n0 101.513
R16272 isrc_sel.n3 isrc_sel 11.8005
R16273 isrc_sel.n3 isrc_sel.n2 4.96991
R16274 isrc_sel.n2 isrc_sel 3.46403
R16275 isrc_sel isrc_sel.n3 2.71109
R16276 vtrip_decoded[0].n0 vtrip_decoded[0].t1 186.374
R16277 vtrip_decoded[0].n0 vtrip_decoded[0].t0 170.308
R16278 vtrip_decoded[0] vtrip_decoded[0].n1 154.56
R16279 vtrip_decoded[0].n2 vtrip_decoded[0].n1 153.462
R16280 vtrip_decoded[0].n1 vtrip_decoded[0].n0 101.513
R16281 vtrip_decoded[0].n3 vtrip_decoded[0] 11.8005
R16282 vtrip_decoded[0].n3 vtrip_decoded[0].n2 4.96991
R16283 vtrip_decoded[0].n2 vtrip_decoded[0] 3.46403
R16284 vtrip_decoded[0] vtrip_decoded[0].n3 2.71109
R16285 vtrip_decoded[5].n0 vtrip_decoded[5].t1 186.374
R16286 vtrip_decoded[5].n0 vtrip_decoded[5].t0 170.308
R16287 vtrip_decoded[5] vtrip_decoded[5].n1 154.56
R16288 vtrip_decoded[5].n2 vtrip_decoded[5].n1 153.462
R16289 vtrip_decoded[5].n1 vtrip_decoded[5].n0 101.513
R16290 vtrip_decoded[5].n3 vtrip_decoded[5] 11.8005
R16291 vtrip_decoded[5].n3 vtrip_decoded[5].n2 4.96991
R16292 vtrip_decoded[5].n2 vtrip_decoded[5] 3.46403
R16293 vtrip_decoded[5] vtrip_decoded[5].n3 2.71109
R16294 vtrip_decoded[7].n0 vtrip_decoded[7].t1 186.374
R16295 vtrip_decoded[7].n0 vtrip_decoded[7].t0 170.308
R16296 vtrip_decoded[7] vtrip_decoded[7].n1 154.56
R16297 vtrip_decoded[7].n2 vtrip_decoded[7].n1 153.462
R16298 vtrip_decoded[7].n1 vtrip_decoded[7].n0 101.513
R16299 vtrip_decoded[7].n3 vtrip_decoded[7] 11.8005
R16300 vtrip_decoded[7].n3 vtrip_decoded[7].n2 4.96991
R16301 vtrip_decoded[7].n2 vtrip_decoded[7] 3.46403
R16302 vtrip_decoded[7] vtrip_decoded[7].n3 2.71109
R16303 ena.n0 ena.t1 186.374
R16304 ena.n0 ena.t0 170.308
R16305 ena ena.n1 154.56
R16306 ena.n2 ena.n1 153.462
R16307 ena.n1 ena.n0 101.513
R16308 ena.n3 ena 11.8005
R16309 ena.n3 ena.n2 4.96991
R16310 ena.n2 ena 3.46403
R16311 ena ena.n3 2.71109
R16312 vtrip_decoded[4].n0 vtrip_decoded[4].t1 186.374
R16313 vtrip_decoded[4].n0 vtrip_decoded[4].t0 170.308
R16314 vtrip_decoded[4] vtrip_decoded[4].n1 154.56
R16315 vtrip_decoded[4].n2 vtrip_decoded[4].n1 153.462
R16316 vtrip_decoded[4].n1 vtrip_decoded[4].n0 101.513
R16317 vtrip_decoded[4].n3 vtrip_decoded[4] 11.8005
R16318 vtrip_decoded[4].n3 vtrip_decoded[4].n2 4.96991
R16319 vtrip_decoded[4].n2 vtrip_decoded[4] 3.46403
R16320 vtrip_decoded[4] vtrip_decoded[4].n3 2.71109
R16321 otrip_decoded[7].n0 otrip_decoded[7].t1 186.374
R16322 otrip_decoded[7].n0 otrip_decoded[7].t0 170.308
R16323 otrip_decoded[7] otrip_decoded[7].n1 154.56
R16324 otrip_decoded[7].n2 otrip_decoded[7].n1 153.462
R16325 otrip_decoded[7].n1 otrip_decoded[7].n0 101.513
R16326 otrip_decoded[7].n3 otrip_decoded[7] 11.8005
R16327 otrip_decoded[7].n3 otrip_decoded[7].n2 4.96991
R16328 otrip_decoded[7].n2 otrip_decoded[7] 3.46403
R16329 otrip_decoded[7] otrip_decoded[7].n3 2.71109
R16330 vtrip_decoded[6].n0 vtrip_decoded[6].t1 186.374
R16331 vtrip_decoded[6].n0 vtrip_decoded[6].t0 170.308
R16332 vtrip_decoded[6] vtrip_decoded[6].n1 154.56
R16333 vtrip_decoded[6].n2 vtrip_decoded[6].n1 153.462
R16334 vtrip_decoded[6].n1 vtrip_decoded[6].n0 101.513
R16335 vtrip_decoded[6].n3 vtrip_decoded[6] 11.8066
R16336 vtrip_decoded[6].n3 vtrip_decoded[6].n2 4.96991
R16337 vtrip_decoded[6].n2 vtrip_decoded[6] 3.46403
R16338 vtrip_decoded[6] vtrip_decoded[6].n3 2.71109
R16339 otrip_decoded[5].n0 otrip_decoded[5].t1 186.374
R16340 otrip_decoded[5].n0 otrip_decoded[5].t0 170.308
R16341 otrip_decoded[5] otrip_decoded[5].n1 154.56
R16342 otrip_decoded[5].n2 otrip_decoded[5].n1 153.462
R16343 otrip_decoded[5].n1 otrip_decoded[5].n0 101.513
R16344 otrip_decoded[5].n3 otrip_decoded[5] 11.8005
R16345 otrip_decoded[5].n3 otrip_decoded[5].n2 4.96991
R16346 otrip_decoded[5].n2 otrip_decoded[5] 3.46403
R16347 otrip_decoded[5] otrip_decoded[5].n3 2.71109
R16348 otrip_decoded[3].n0 otrip_decoded[3].t1 186.374
R16349 otrip_decoded[3].n0 otrip_decoded[3].t0 170.308
R16350 otrip_decoded[3] otrip_decoded[3].n1 154.56
R16351 otrip_decoded[3].n2 otrip_decoded[3].n1 153.462
R16352 otrip_decoded[3].n1 otrip_decoded[3].n0 101.513
R16353 otrip_decoded[3].n3 otrip_decoded[3] 11.8005
R16354 otrip_decoded[3].n3 otrip_decoded[3].n2 4.96991
R16355 otrip_decoded[3].n2 otrip_decoded[3] 3.46403
R16356 otrip_decoded[3] otrip_decoded[3].n3 2.71109
R16357 otrip_decoded[1].n0 otrip_decoded[1].t1 186.374
R16358 otrip_decoded[1].n0 otrip_decoded[1].t0 170.308
R16359 otrip_decoded[1] otrip_decoded[1].n1 154.56
R16360 otrip_decoded[1].n2 otrip_decoded[1].n1 153.462
R16361 otrip_decoded[1].n1 otrip_decoded[1].n0 101.513
R16362 otrip_decoded[1].n3 otrip_decoded[1] 11.8005
R16363 otrip_decoded[1].n3 otrip_decoded[1].n2 4.96991
R16364 otrip_decoded[1].n2 otrip_decoded[1] 3.46403
R16365 otrip_decoded[1] otrip_decoded[1].n3 2.71109
C0 rstring_mux_0.otrip_decoded_b_avdd[2] avss 0.363375f
C1 a_n13099_n19314# avss 0.466333f
C2 rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.otrip_decoded_b_avdd[3] 0.155509f
C3 a_n11975_9395# a_n11219_9395# 0.296258f
C4 a_n1783_n2964# a_n1683_n2876# 0.40546f
C5 comparator_0.ena a_10084_n3212# 0.137017f
C6 rc_osc_0.in rc_osc_0.m 1.10731f
C7 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_avdd[4] 0.503487f
C8 ibias_gen_0.ena_b ibg_200n 0.467695f
C9 a_n3527_n3946# dvdd 0.176016f
C10 ibias_gen_0.ibias0 avss 1.14866f
C11 a_8777_n2964# dvdd 0.380862f
C12 a_n10075_n19314# a_n9319_n19314# 0.296258f
C13 rstring_mux_0.otrip_decoded_avdd[1] avss 1.63066f
C14 rstring_mux_0.otrip_decoded_b_avdd[3] avdd 0.903548f
C15 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip2 0.190544f
C16 rstring_mux_0.otrip_decoded_avdd[3] avdd 1.72135f
C17 a_2399_n11914# a_3155_n11914# 0.296258f
C18 a_n5161_n11914# vin_vunder 0.159467f
C19 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[2] 0.10426f
C20 a_1636_n3212# rstring_mux_0.vtrip_decoded_avdd[0] 0.135959f
C21 a_n8119_n1230# otrip_decoded[1] 0.207169f
C22 a_n1415_n3946# avdd 0.143952f
C23 rstring_mux_0.vtrip4 avss 2.05606f
C24 comparator_0.ena ibias_gen_0.vp1 0.338208f
C25 rstring_mux_0.vtrip2 vin_vunder 2.31192f
C26 a_8877_n2876# avdd 0.864301f
C27 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X rstring_mux_0.otrip_decoded_avdd[3] 1.37931f
C28 rstring_mux_0.otrip_decoded_avdd[2] dvdd 0.255576f
C29 a_4921_n2212# dvdd 0.169343f
C30 a_n1783_n2964# a_n1415_n3946# 0.138963f
C31 a_n1783_n1230# a_n1683_n1142# 0.40546f
C32 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip_decoded_b_avdd[4] 0.154961f
C33 a_n10453_n11914# vin_vunder 0.159467f
C34 rstring_mux_0.vtrip_decoded_avdd[1] dcomp3v3uv 0.100293f
C35 rstring_mux_0.otrip_decoded_b_avdd[2] vin_brout 0.34139f
C36 a_1636_n1478# rstring_mux_0.vtrip_decoded_avdd[1] 0.13699f
C37 a_n476_n1478# avdd 0.420074f
C38 a_n15367_n19314# a_n14611_n19314# 0.296258f
C39 dcomp3v3uv avss 7.27403f
C40 a_11121_n23089# a_11121_n23845# 0.296258f
C41 vl schmitt_trigger_0.in 0.503663f
C42 a_n4405_n11914# a_n3649_n11914# 0.296258f
C43 a_n15745_n11914# vin_vunder 0.161624f
C44 ibias_gen_0.ibias0 vin_brout 2.74533f
C45 rstring_mux_0.otrip_decoded_avdd[1] vin_brout 0.881159f
C46 a_7691_n11914# avss 0.525451f
C47 a_n22294_n2937# avss 0.471605f
C48 ibias_gen_0.isrc_sel dvdd 0.176564f
C49 a_7458_n3990# a_7033_n3946# 0.460766f
C50 comparator_0.ena ibias_gen_0.ibias0 1.70445f
C51 comparator_0.ena rstring_mux_0.otrip_decoded_avdd[1] 0.17335f
C52 ibias_gen_0.isrc_sel_b avdd 3.36468f
C53 vl dvdd 1.96235f
C54 rstring_mux_0.vtrip_decoded_b_avdd[6] vin_vunder 0.340862f
C55 a_8777_n2964# a_8877_n2876# 0.40546f
C56 rstring_mux_0.vtrip4 vin_brout 2.26482f
C57 a_n9329_1995# a_n8573_1995# 0.296258f
C58 rstring_mux_0.vtop a_n15745_n11914# 0.348335f
C59 a_n11975_9395# avss 0.460203f
C60 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_avdd[2] 1.42613f
C61 a_329_n2964# avdd 0.207177f
C62 a_n24940_n10337# a_n24184_n10337# 0.296258f
C63 comparator_0.n0 vbg_1v2 0.692613f
C64 a_2399_n11914# avss 0.465592f
C65 comparator_1.vpp comparator_1.vn 0.327643f
C66 comparator_1.ena_b avdd 0.998725f
C67 a_5045_n19314# a_5801_n19314# 0.296258f
C68 ibias_gen_0.ena_b ibias_gen_0.isrc_sel 1.07804f
C69 a_10084_n1478# avdd 0.418567f
C70 a_n1683_n2876# a_n476_n3212# 0.28899f
C71 rstring_mux_0.otrip_decoded_b_avdd[7] avss 0.36282f
C72 a_697_n3946# dvdd 0.176016f
C73 rc_osc_0.vr osc_ena 0.245726f
C74 a_n3895_n2964# otrip_decoded[4] 0.2082f
C75 rstring_mux_0.vtrip_decoded_avdd[7] avss 1.38048f
C76 a_n9697_n11914# a_n8941_n11914# 0.296258f
C77 a_5346_n2256# avdd 0.607928f
C78 a_n4405_n11914# avss 0.482553f
C79 a_8777_n1230# isrc_sel 0.2082f
C80 a_8777_n1230# a_8877_n1142# 0.40546f
C81 avdd vbg_1v2 8.1878f
C82 rstring_mux_0.vtrip_decoded_b_avdd[0] avdd 0.903548f
C83 comparator_0.ena dcomp3v3uv 0.508881f
C84 a_2809_n3946# avdd 0.143952f
C85 a_n9329_1995# avss 0.460231f
C86 rstring_mux_0.vtrip6 avss 2.27146f
C87 rstring_mux_0.vtrip4 vin_vunder 2.34032f
C88 a_n14621_1995# a_n13865_1995# 0.296258f
C89 rstring_mux_0.otrip_decoded_avdd[0] avdd 1.34894f
C90 comparator_1.vn avss 8.76998f
C91 a_n24940_n10337# avss 0.472978f
C92 a_5346_n3990# dvdd 0.104499f
C93 a_5045_n19314# avss 0.466333f
C94 a_7033_n2212# dvdd 0.169343f
C95 rc_osc_0.in rc_osc_0.vr 0.495731f
C96 a_n1683_n1142# a_n476_n1478# 0.28899f
C97 a_n9697_n11914# avss 0.465068f
C98 rstring_mux_0.vtrip_decoded_avdd[4] rstring_mux_0.vtrip_decoded_b_avdd[3] 0.155115f
C99 a_n247_n19314# a_509_n19314# 0.296258f
C100 a_329_n1230# dvdd 0.379209f
C101 a_10514_n2760# avdd 0.53813f
C102 a_n14621_1995# avss 0.4604f
C103 a_9145_n2212# avdd 0.143323f
C104 a_n247_n19314# avss 0.466333f
C105 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip0 0.190544f
C106 ibias_gen_0.vp1 ibias_gen_0.ena_b 0.142844f
C107 a_429_n1142# avdd 0.863296f
C108 a_n14989_n11914# a_n14233_n11914# 0.296258f
C109 a_5860_n3212# rstring_mux_0.vtrip_decoded_avdd[4] 0.135915f
C110 rstring_mux_0.otrip_decoded_avdd[0] rstring_mux_0.vtrip0 0.50883f
C111 a_n14989_n11914# avss 0.465096f
C112 a_n10279_n23467# a_n10279_n24223# 0.296258f
C113 rstring_mux_0.otrip_decoded_b_avdd[7] vin_brout 0.340862f
C114 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[1] 0.556851f
C115 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_b_avdd[7] 0.572384f
C116 a_9570_n3990# a_9145_n3946# 0.460766f
C117 comparator_0.ena rstring_mux_0.vtrip_decoded_avdd[7] 1.91505f
C118 a_n16775_n2223# avdd 0.466408f
C119 a_6665_n2964# a_7033_n3946# 0.138963f
C120 rc_osc_0.ena_b dvdd 0.500996f
C121 a_n7051_n19314# avss 0.466333f
C122 rstring_mux_0.otrip_decoded_avdd[1] dvdd 0.266224f
C123 a_8877_n2876# a_10084_n3212# 0.28899f
C124 rstring_mux_0.vtrip6 vin_brout 2.08469f
C125 a_n8951_9395# a_n8195_9395# 0.296258f
C126 a_n7051_n19314# a_n6295_n19314# 0.296258f
C127 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b 1.79811f
C128 comparator_0.vt comparator_0.vnn 4.29222f
C129 rstring_mux_0.vtrip_decoded_avdd[5] avss 1.50537f
C130 a_5346_n2256# a_4921_n2212# 0.460766f
C131 a_1636_n3212# avdd 0.421965f
C132 rc_osc_0.in avdd 0.210176f
C133 a_n24562_n2937# a_n23806_n2937# 0.296258f
C134 comparator_1.n0 dcomp3v3 0.945307f
C135 comparator_0.ena comparator_1.vn 0.293425f
C136 comparator_1.vpp comparator_1.n0 0.347877f
C137 comparator_1.vnn comparator_1.vm 0.563119f
C138 a_5423_n11914# a_6179_n11914# 0.296258f
C139 comparator_1.vt dcomp3v3 2.36366f
C140 comparator_1.vt comparator_1.vpp 2.58192f
C141 a_3234_n2256# avdd 0.607928f
C142 a_5860_n1478# rstring_mux_0.vtrip_decoded_avdd[5] 0.13699f
C143 a_n6007_n1230# a_n5639_n2212# 0.138963f
C144 a_n12343_n19314# avss 0.466333f
C145 rstring_mux_0.otrip_decoded_avdd[5] dcomp3v3uv 0.213252f
C146 ibias_gen_0.isrc_sel a_10084_n1478# 0.155566f
C147 a_4921_n3946# dvdd 0.176016f
C148 a_n6007_n1230# otrip_decoded[3] 0.207704f
C149 a_3234_n3990# dvdd 0.104499f
C150 rstring_mux_0.vtrip_decoded_avdd[7] vin_vunder 0.880681f
C151 a_10874_n1026# avdd 0.177477f
C152 a_8877_n1142# a_10084_n1478# 0.28899f
C153 a_n4405_n11914# vin_vunder 0.157512f
C154 rstring_mux_0.vtrip_decoded_b_avdd[4] avss 0.36282f
C155 schmitt_trigger_0.in dcomp3v3uv 0.122613f
C156 dcomp3v3uv comparator_0.n1 1.71428f
C157 a_n8119_n1230# avdd 0.194982f
C158 sky130_fd_sc_hd__inv_4_3.Y dcomp 1.48254f
C159 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_b_avdd[2] 0.155546f
C160 comparator_0.vpp avss 2.27913f
C161 rstring_mux_0.vtrip_decoded_avdd[6] avdd 1.9364f
C162 rstring_mux_0.vtrip6 vin_vunder 2.27059f
C163 a_n14243_9395# a_n13487_9395# 0.296258f
C164 comparator_1.n0 avss 3.94229f
C165 dcomp3v3uv dvdd 1.09406f
C166 comparator_1.vt avss 29.094501f
C167 rstring_mux_0.vtrip_decoded_b_avdd[5] avdd 0.90363f
C168 a_n12343_n19314# a_n11587_n19314# 0.296258f
C169 a_6765_n1142# a_7458_n2256# 0.264594f
C170 a_n8119_n2964# dvdd 0.382499f
C171 a_329_n2964# a_697_n3946# 0.138963f
C172 rstring_mux_0.otrip_decoded_b_avdd[0] avss 0.399825f
C173 a_131_n11914# a_887_n11914# 0.296258f
C174 a_n9697_n11914# vin_vunder 0.128847f
C175 ibias_gen_0.vp1 ibias_gen_0.isrc_sel_b 0.406323f
C176 a_n8019_n2876# avdd 0.864385f
C177 a_1122_n2256# a_697_n2212# 0.460766f
C178 rstring_mux_0.otrip_decoded_b_avdd[1] avdd 0.904297f
C179 a_2441_n1230# avdd 0.206171f
C180 a_n5907_n2876# a_n5214_n3990# 0.264594f
C181 a_n14989_n11914# vin_vunder 0.159695f
C182 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[7] 0.377385f
C183 comparator_0.ibias a_n26830_n2937# 0.134538f
C184 a_n21916_n10337# a_n21160_n10337# 0.296258f
C185 a_n21538_n2937# avss 0.471774f
C186 a_8447_n11914# avss 0.525755f
C187 a_8069_n19314# a_8825_n19314# 0.296258f
C188 rstring_mux_0.vtrip_decoded_avdd[3] avss 1.48249f
C189 dvdd vunder 1.54357f
C190 rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.otrip_decoded_b_avdd[6] 0.573474f
C191 a_1122_n2256# avdd 0.607928f
C192 a_2441_n2964# dvdd 0.380879f
C193 rstring_mux_0.vtrip_decoded_avdd[7] dvdd 0.289581f
C194 comparator_0.vpp comparator_0.vm 0.636921f
C195 comparator_0.vnn comparator_0.vn 0.298803f
C196 rstring_mux_0.otrip_decoded_avdd[3] dcomp3v3uv 0.156703f
C197 a_n6673_n11914# a_n5917_n11914# 0.296258f
C198 comparator_1.vt vin_brout 25.678198f
C199 a_n11219_9395# avss 0.460203f
C200 ibias_gen_0.isrc_sel a_n16775_n2223# 0.291728f
C201 comparator_0.vt comparator_0.vn 0.209988f
C202 comparator_0.ena comparator_0.vpp 0.609928f
C203 a_10515_n1026# a_10515_n2156# 0.170258f
C204 a_2541_n2876# avdd 0.863791f
C205 a_1122_n3990# dvdd 0.104499f
C206 a_3155_n11914# avss 0.465978f
C207 rstring_mux_0.vtrip_decoded_avdd[5] vin_vunder 0.878049f
C208 comparator_0.ena comparator_1.n0 0.123113f
C209 a_n26830_n2937# avss 0.776278f
C210 comparator_1.vt comparator_0.ena 0.306818f
C211 rstring_mux_0.otrip_decoded_b_avdd[0] vin_brout 0.343304f
C212 a_7458_n2256# dvdd 0.104499f
C213 a_n15529_n2223# ibg_200n 0.397003f
C214 a_n5907_n1142# a_n5214_n2256# 0.264594f
C215 comparator_0.ibias itest 0.10252f
C216 a_n1783_n2964# otrip_decoded[6] 0.2082f
C217 comparator_0.ibias comparator_0.ena_b 0.195795f
C218 a_329_n2964# a_429_n2876# 0.40546f
C219 a_n11597_1995# a_n10841_1995# 0.296258f
C220 rstring_mux_0.vtrip_decoded_avdd[4] avdd 1.61396f
C221 a_7033_n3946# dvdd 0.176016f
C222 a_n9697_n11914# dvdd 0.431259f
C223 rstring_mux_0.vtrip_decoded_avdd[7] rstring_mux_0.vtrip_decoded_b_avdd[7] 0.572453f
C224 a_n3102_n2256# a_n3527_n2212# 0.460766f
C225 comparator_1.ena_b ibias_gen_0.ibias0 0.201284f
C226 a_9570_n2256# avdd 0.612302f
C227 comparator_1.vm avdd 0.382522f
C228 a_n27208_n10337# a_n26452_n10337# 0.296258f
C229 a_n3649_n11914# avss 0.465525f
C230 a_2777_n19314# a_3533_n19314# 0.296258f
C231 rstring_mux_0.vtrip_decoded_b_avdd[4] vin_vunder 0.340862f
C232 a_n6812_n1478# avdd 0.420451f
C233 a_9145_n3946# avdd 0.144336f
C234 a_n8573_1995# avss 0.4604f
C235 rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.otrip_decoded_b_avdd[1] 0.155388f
C236 comparator_0.ena_b avss 1.76426f
C237 comparator_0.vpp vin_vunder 2.49904f
C238 a_n24184_n10337# avss 0.472978f
C239 dcomp3v3 avss 3.78523f
C240 comparator_1.vpp avss 1.79171f
C241 a_5801_n19314# avss 0.466333f
C242 a_n11965_n11914# a_n11209_n11914# 0.296258f
C243 a_329_n1230# a_429_n1142# 0.40546f
C244 a_n8941_n11914# avss 0.465068f
C245 comparator_0.ibias avss 4.73461f
C246 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[5] 0.174324f
C247 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_avdd[0] 3.24722f
C248 a_n13865_1995# avss 0.460231f
C249 a_n14999_9395# a_n14243_9395# 0.296258f
C250 rstring_mux_0.otrip_decoded_b_avdd[5] avss 0.36282f
C251 a_n6007_n2964# avdd 0.207177f
C252 rstring_mux_0.vtrip_decoded_avdd[1] avss 1.39274f
C253 a_509_n19314# avss 0.466333f
C254 a_n990_n2256# avdd 0.607928f
C255 a_3748_n1478# avdd 0.420074f
C256 rstring_mux_0.vtrip_decoded_avdd[5] dvdd 0.324294f
C257 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip_decoded_b_avdd[2] 0.155157f
C258 rstring_mux_0.otrip_decoded_b_avdd[6] avdd 0.903548f
C259 a_n14233_n11914# avss 0.465264f
C260 a_n21538_n2937# a_n20782_n2937# 0.296258f
C261 a_8447_n11914# a_9203_n11914# 0.296258f
C262 a_n990_n3990# dvdd 0.104499f
C263 a_n7326_n2256# a_n7751_n2212# 0.460766f
C264 rstring_mux_0.vtrip_decoded_avdd[3] vin_vunder 0.879435f
C265 a_3234_n3990# a_2809_n3946# 0.460766f
C266 a_8777_n2964# a_9145_n3946# 0.138963f
C267 a_n6295_n19314# avss 0.466333f
C268 rc_osc_0.ena_b osc_ena 0.488092f
C269 comparator_0.vnn comparator_0.n0 0.428003f
C270 dvdd outb 1.54606f
C271 schmitt_trigger_0.in comparator_0.vpp 0.250959f
C272 a_10873_n2760# avdd 0.177483f
C273 comparator_0.ena comparator_0.ena_b 0.623387f
C274 rstring_mux_0.vtrip_decoded_avdd[2] avdd 1.66091f
C275 comparator_1.vpp vin_brout 2.54645f
C276 comparator_0.ena itest 0.154848f
C277 dcomp3v3uv vbg_1v2 0.3098f
C278 a_4553_n2964# avdd 0.207177f
C279 comparator_1.vpp comparator_0.ena 0.784496f
C280 a_n3895_n1230# a_n3527_n2212# 0.138963f
C281 rc_osc_0.m rc_osc_0.vr 0.559422f
C282 dvdd osc_ck 1.35201f
C283 a_10874_n2222# dvdd 0.469294f
C284 a_n3895_n1230# otrip_decoded[5] 0.2082f
C285 a_n1683_n2876# a_n990_n3990# 0.264594f
C286 a_n11587_n19314# avss 0.466333f
C287 a_n6007_n1230# dvdd 0.385817f
C288 a_429_n2876# a_1636_n3212# 0.28899f
C289 a_n11219_9395# a_n10463_9395# 0.296258f
C290 rstring_mux_0.otrip_decoded_b_avdd[5] vin_brout 0.340862f
C291 comparator_0.ena comparator_0.ibias 3.0153f
C292 rc_osc_0.ena_b rc_osc_0.in 0.13356f
C293 comparator_0.vnn avdd 37.3266f
C294 a_n9319_n19314# a_n8563_n19314# 0.296258f
C295 rstring_mux_0.vtrip_decoded_avdd[6] rstring_mux_0.vtrip_decoded_b_avdd[6] 0.572868f
C296 sky130_fd_sc_hd__inv_4_1.Y vunder 1.48088f
C297 comparator_1.n1 avdd 2.69603f
C298 a_n7751_n2212# avdd 0.142924f
C299 a_10514_n2760# dcomp3v3uv 0.223996f
C300 comparator_0.vt avdd 0.142093p
C301 a_n26830_n2937# a_n26074_n2937# 0.296258f
C302 a_3155_n11914# a_3911_n11914# 0.296258f
C303 a_n3649_n11914# vin_vunder 0.154012f
C304 a_n5907_n1142# avdd 0.863296f
C305 avss vin_brout 14.4003f
C306 comparator_0.vm avss 10.3984f
C307 vl sky130_fd_sc_hd__inv_4_3.Y 0.396105f
C308 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[3] 0.14576f
C309 comparator_0.ena avss 19.7509f
C310 rstring_mux_0.otrip_decoded_avdd[7] avss 1.37218f
C311 comparator_1.ena_b comparator_1.vn 1.12092f
C312 rstring_mux_0.vtrip0 a_n4027_n19314# 0.298434f
C313 a_8877_n1142# a_9570_n2256# 0.264594f
C314 a_n990_n3990# a_n1415_n3946# 0.460766f
C315 a_n3102_n2256# avdd 0.607928f
C316 a_n1683_n1142# a_n990_n2256# 0.264594f
C317 a_2441_n2964# a_2809_n3946# 0.138963f
C318 rstring_mux_0.vtrip_decoded_avdd[3] dvdd 0.517826f
C319 a_429_n1142# a_1636_n1478# 0.28899f
C320 a_n8941_n11914# vin_vunder 0.128847f
C321 a_4553_n1230# dvdd 0.379209f
C322 a_n4700_n3212# avdd 0.421965f
C323 a_10515_n1026# a_10874_n1026# 0.249533f
C324 a_n3102_n3990# dvdd 0.104499f
C325 rstring_mux_0.vtrip_decoded_avdd[1] vin_vunder 0.909999f
C326 comparator_1.vn vbg_1v2 0.723918f
C327 a_n14611_n19314# a_n13855_n19314# 0.296258f
C328 a_4653_n1142# avdd 0.863296f
C329 rstring_mux_0.vtrip_decoded_b_avdd[2] avss 0.362817f
C330 rstring_mux_0.vtrip_decoded_avdd[2] rstring_mux_0.vtrip_decoded_b_avdd[1] 0.155018f
C331 a_11121_n23845# a_11121_n24601# 0.296258f
C332 a_n14233_n11914# vin_vunder 0.159467f
C333 a_n20782_n2937# avss 0.47927f
C334 rstring_mux_0.vtrip_decoded_avdd[0] avdd 1.59456f
C335 a_9203_n11914# avss 0.82426f
C336 a_7458_n3990# dvdd 0.104499f
C337 avss vin_vunder 10.8061f
C338 rstring_mux_0.vtrip_decoded_b_avdd[3] avdd 0.903548f
C339 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_b_avdd[1] 0.569059f
C340 comparator_0.vn comparator_0.n0 1.99139f
C341 a_n8573_1995# schmitt_trigger_0.in 0.303942f
C342 a_9570_n3990# avdd 0.61228f
C343 rstring_mux_0.vtop avss 3.67651f
C344 comparator_0.ena vin_brout 2.34883f
C345 a_n10463_9395# avss 0.460203f
C346 rstring_mux_0.otrip_decoded_avdd[7] vin_brout 0.875535f
C347 a_5860_n3212# avdd 0.421965f
C348 a_10874_n2222# a_10515_n2156# 0.249269f
C349 a_329_n2964# vtrip_decoded[0] 0.2082f
C350 a_n26074_n2937# avss 0.484544f
C351 a_n24184_n10337# a_n23428_n10337# 0.296258f
C352 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_b_avdd[5] 0.573322f
C353 a_5801_n19314# a_6557_n19314# 0.296258f
C354 a_3911_n11914# avss 0.484363f
C355 rstring_mux_0.vtrip_decoded_avdd[6] dcomp3v3uv 0.194356f
C356 a_n5214_n3990# a_n5639_n3946# 0.460766f
C357 a_n5639_n2212# dvdd 0.16995f
C358 dcomp3v3 dvdd 1.10728f
C359 rstring_mux_0.vtrip_decoded_avdd[0] rstring_mux_0.vtrip0 0.485675f
C360 schmitt_trigger_0.in schmitt_trigger_0.m 0.957373f
C361 a_n6812_n3212# rstring_mux_0.otrip_decoded_avdd[0] 0.135767f
C362 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[1] 0.133642f
C363 comparator_0.vn avdd 0.753795f
C364 a_n8941_n11914# a_n8185_n11914# 0.296258f
C365 rstring_mux_0.otrip_decoded_avdd[5] avss 1.34873f
C366 a_n3527_n2212# avdd 0.142934f
C367 schmitt_trigger_0.m dvdd 2.69554f
C368 comparator_1.vnn avdd 37.3119f
C369 a_n5214_n2256# avdd 0.607928f
C370 a_n3895_n1230# avdd 0.206171f
C371 rstring_mux_0.vtrip_decoded_avdd[1] dvdd 0.335417f
C372 rstring_mux_0.vtrip_decoded_avdd[2] rstring_mux_0.vtrip2 0.4803f
C373 a_n4700_n3212# rstring_mux_0.otrip_decoded_avdd[2] 0.135981f
C374 schmitt_trigger_0.in avss 8.82092f
C375 comparator_0.n1 avss 3.03066f
C376 vin_brout vin_vunder 0.868683f
C377 a_n8119_n2964# a_n8019_n2876# 0.40546f
C378 a_n13865_1995# a_n13109_1995# 0.296258f
C379 a_n23428_n10337# avss 0.472978f
C380 a_n5214_n3990# dvdd 0.104499f
C381 a_6557_n19314# avss 0.466333f
C382 comparator_0.ena vin_vunder 0.229267f
C383 ibias_gen_0.ibias0 comparator_1.vm 0.155341f
C384 a_n3895_n2964# dvdd 0.380879f
C385 avss dvdd 2.52914f
C386 a_n8185_n11914# avss 0.465068f
C387 a_509_n19314# a_1265_n19314# 0.296258f
C388 a_2541_n2876# a_3234_n3990# 0.264594f
C389 a_n6812_n1478# rstring_mux_0.otrip_decoded_avdd[1] 0.13699f
C390 rstring_mux_0.vtrip_decoded_avdd[4] rstring_mux_0.vtrip4 0.497379f
C391 rstring_mux_0.vtrip_decoded_avdd[7] rstring_mux_0.vtrip_decoded_avdd[6] 3.06282f
C392 rstring_mux_0.otrip_decoded_avdd[6] avdd 1.62903f
C393 a_n13109_1995# avss 0.460203f
C394 a_n3795_n2876# avdd 0.863791f
C395 comparator_0.vpp vbg_1v2 2.95415f
C396 a_1265_n19314# avss 0.466333f
C397 comparator_1.n0 vbg_1v2 0.530131f
C398 a_n14233_n11914# a_n13477_n11914# 0.296258f
C399 a_6665_n1230# avdd 0.206171f
C400 comparator_1.vt vbg_1v2 24.6722f
C401 rstring_mux_0.vtrip_decoded_b_avdd[2] vin_vunder 0.340862f
C402 rstring_mux_0.vtrip_decoded_avdd[6] rstring_mux_0.vtrip6 0.488466f
C403 a_n4700_n1478# rstring_mux_0.otrip_decoded_avdd[3] 0.13699f
C404 a_n13477_n11914# avss 0.466481f
C405 a_n8119_n1230# a_n8019_n1142# 0.40546f
C406 ibias_gen_0.ena_b avss 2.71238f
C407 a_n10279_n24223# a_n10279_n24979# 0.296258f
C408 rstring_mux_0.vtrip_decoded_b_avdd[7] avss 0.479446f
C409 rstring_mux_0.otrip_decoded_avdd[5] vin_brout 0.876971f
C410 a_10873_n3956# dvdd 0.469495f
C411 a_6665_n2964# dvdd 0.380879f
C412 a_2541_n1142# a_3234_n2256# 0.264594f
C413 rstring_mux_0.vtrip_decoded_avdd[4] dcomp3v3uv 0.249577f
C414 rstring_mux_0.otrip_decoded_avdd[0] rstring_mux_0.otrip_decoded_b_avdd[0] 0.56463f
C415 a_n5539_n19314# avss 0.466333f
C416 rstring_mux_0.ena_b avdd 6.38079f
C417 a_n7751_n3946# avdd 0.143941f
C418 a_n6295_n19314# a_n5539_n19314# 0.296258f
C419 comparator_0.ena schmitt_trigger_0.in 1.21644f
C420 rstring_mux_0.vtop vin_vunder 1.24609f
C421 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[7] 0.126209f
C422 a_n1783_n1230# otrip_decoded[7] 0.2082f
C423 rstring_mux_0.otrip_decoded_b_avdd[3] avss 0.362817f
C424 a_6765_n2876# avdd 0.863791f
C425 a_n23806_n2937# a_n23050_n2937# 0.296258f
C426 a_6179_n11914# a_6935_n11914# 0.296258f
C427 rstring_mux_0.otrip_decoded_avdd[3] avss 1.341f
C428 dvdd vin_brout 0.119455f
C429 rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.otrip_decoded_b_avdd[4] 0.57199f
C430 a_n1783_n1230# a_n1415_n2212# 0.138963f
C431 a_n1415_n2212# dvdd 0.169343f
C432 a_n7326_n2256# avdd 0.607831f
C433 comparator_0.ena dvdd 0.351058f
C434 rstring_mux_0.otrip_decoded_avdd[7] dvdd 0.291769f
C435 a_n10831_n19314# avss 0.466333f
C436 osc_ena osc_ck 0.143345f
C437 rstring_mux_0.otrip_decoded_b_avdd[4] avdd 0.903548f
C438 a_2441_n2964# a_2541_n2876# 0.40546f
C439 comparator_0.n0 avdd 1.07016f
C440 a_n7326_n3990# dvdd 0.104499f
C441 sky130_fd_sc_hd__inv_4_4.Y outb 1.48254f
C442 a_697_n2212# avdd 0.142934f
C443 a_n2588_n1478# avdd 0.420074f
C444 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip_decoded_avdd[6] 1.33995f
C445 a_n16123_n19314# avss 0.732759f
C446 comparator_0.ena ibias_gen_0.ena_b 1.24167f
C447 a_n8019_n2876# a_n6812_n3212# 0.28899f
C448 rstring_mux_0.otrip_decoded_avdd[4] avdd 1.52975f
C449 a_n13487_9395# a_n12731_9395# 0.296258f
C450 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip_decoded_b_avdd[5] 0.574941f
C451 rc_osc_0.in osc_ck 1.05774f
C452 comparator_0.ena rstring_mux_0.vtrip_decoded_b_avdd[7] 0.1256f
C453 a_n11587_n19314# a_n10831_n19314# 0.296258f
C454 a_4553_n2964# a_4921_n3946# 0.138963f
C455 dvdd vin_vunder 0.119455f
C456 a_2441_n1230# a_2541_n1142# 0.40546f
C457 a_887_n11914# a_1643_n11914# 0.296258f
C458 a_n8185_n11914# vin_vunder 0.159467f
C459 rstring_mux_0.otrip_decoded_b_avdd[3] vin_brout 0.340862f
C460 rstring_mux_0.otrip_decoded_avdd[3] vin_brout 0.880782f
C461 a_10874_n1026# a_10874_n2222# 0.136815f
C462 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X avdd 3.01562f
C463 a_n1783_n2964# avdd 0.207177f
C464 comparator_1.vn comparator_1.vm 4.6608f
C465 ibias_gen_0.isrc_sel_b avss 2.66768f
C466 rstring_mux_0.vtop dvdd 0.177165f
C467 rstring_mux_0.vtrip_decoded_avdd[2] dcomp3v3uv 0.359441f
C468 comparator_1.vpp vbg_1v2 3.00457f
C469 avdd ibg_200n 0.695438f
C470 a_7972_n1478# avdd 0.420074f
C471 a_n476_n3212# rstring_mux_0.otrip_decoded_avdd[6] 0.136228f
C472 a_n8019_n1142# a_n6812_n1478# 0.28899f
C473 a_n13477_n11914# vin_vunder 0.159467f
C474 a_n21160_n10337# a_n20404_n10337# 0.296258f
C475 rstring_mux_0.vtrip_decoded_b_avdd[7] vin_vunder 0.340862f
C476 a_8825_n19314# a_9581_n19314# 0.296258f
C477 a_n5639_n3946# dvdd 0.176016f
C478 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[5] 0.101776f
C479 rstring_mux_0.vtrip0 avdd 0.430845f
C480 comparator_1.ena_b avss 1.77799f
C481 a_2441_n2964# vtrip_decoded[2] 0.2082f
C482 rstring_mux_0.otrip_decoded_avdd[5] dvdd 0.42314f
C483 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip_decoded_b_avdd[0] 0.155269f
C484 a_n3527_n3946# avdd 0.143952f
C485 a_n5917_n11914# a_n5161_n11914# 0.296258f
C486 a_n9707_9395# avss 0.460203f
C487 a_8777_n2964# avdd 0.207184f
C488 a_n25318_n2937# avss 0.472952f
C489 schmitt_trigger_0.in dvdd 2.6898f
C490 a_4667_n11914# avss 0.525451f
C491 avss vbg_1v2 11.1373f
C492 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.vtrip6 0.190544f
C493 a_2809_n2212# dvdd 0.169343f
C494 a_n476_n1478# rstring_mux_0.otrip_decoded_avdd[7] 0.13699f
C495 rstring_mux_0.vtrip_decoded_b_avdd[0] avss 0.36282f
C496 a_n1783_n1230# dvdd 0.387197f
C497 a_n10841_1995# a_n10085_1995# 0.296258f
C498 a_2541_n2876# a_3748_n3212# 0.28899f
C499 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip_decoded_avdd[4] 2.29102f
C500 rstring_mux_0.otrip_decoded_avdd[0] avss 1.64125f
C501 rstring_mux_0.otrip_decoded_avdd[2] avdd 1.52848f
C502 rstring_mux_0.vtrip_decoded_b_avdd[1] avdd 0.903548f
C503 a_4921_n2212# avdd 0.142934f
C504 a_n26452_n10337# a_n25696_n10337# 0.296258f
C505 comparator_0.ena ibias_gen_0.isrc_sel_b 1.98919f
C506 a_3533_n19314# a_4289_n19314# 0.296258f
C507 a_n1683_n1142# avdd 0.863296f
C508 sky130_fd_sc_hd__inv_4_1.A dvdd 0.677586f
C509 a_7313_n19314# avss 0.466333f
C510 a_n22672_n10337# avss 0.472978f
C511 comparator_0.ena comparator_1.ena_b 0.706636f
C512 a_6665_n1230# a_7033_n2212# 0.138963f
C513 comparator_1.vnn ibias_gen_0.ibias0 1.84751f
C514 rstring_mux_0.vtrip_decoded_avdd[4] rstring_mux_0.vtrip_decoded_b_avdd[4] 0.572505f
C515 a_n11209_n11914# a_n10453_n11914# 0.296258f
C516 rstring_mux_0.vtrip_decoded_avdd[0] dcomp3v3uv 0.49775f
C517 a_2541_n1142# a_3748_n1478# 0.28899f
C518 a_n7429_n11914# avss 0.465068f
C519 a_8777_n1230# dvdd 0.379192f
C520 ibias_gen_0.isrc_sel avdd 10.4627f
C521 a_n12353_1995# avss 0.460203f
C522 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[3] 0.117015f
C523 a_n476_n3212# avdd 0.421965f
C524 vin_brout vbg_1v2 7.42266f
C525 comparator_1.vm comparator_1.n0 2.59034f
C526 a_2021_n19314# avss 0.466333f
C527 vl avdd 2.35468f
C528 a_10514_n2760# a_10873_n3956# 0.166612f
C529 rc_osc_0.vr a_n10279_n22711# 0.301135f
C530 comparator_0.ena vbg_1v2 0.553802f
C531 a_8877_n1142# avdd 0.863813f
C532 comparator_0.ena rstring_mux_0.vtrip_decoded_b_avdd[0] 0.100519f
C533 rstring_mux_0.otrip_decoded_avdd[3] dvdd 0.382485f
C534 rstring_mux_0.otrip_decoded_avdd[0] vin_brout 0.882514f
C535 a_n12721_n11914# avss 0.466465f
C536 rc_osc_0.in a_n10279_n24223# 0.516433f
C537 vl sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 0.799678f
C538 comparator_0.ena rstring_mux_0.otrip_decoded_avdd[0] 0.826776f
C539 a_n1415_n3946# dvdd 0.176016f
C540 rc_osc_0.in avss 0.362331f
C541 rstring_mux_0.vtrip2 avdd 0.859231f
C542 a_n4783_n19314# avss 0.466333f
C543 a_329_n1230# vtrip_decoded[1] 0.2082f
C544 dvdd brout_filt 1.55425f
C545 rstring_mux_0.vtrip_decoded_avdd[0] rstring_mux_0.otrip_decoded_b_avdd[7] 0.154952f
C546 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip_decoded_avdd[4] 1.04751f
C547 a_697_n3946# avdd 0.143952f
C548 a_10084_n3212# avdd 0.420425f
C549 a_329_n1230# a_697_n2212# 0.138963f
C550 vbg_1v2 vin_vunder 4.30452f
C551 rc_osc_0.ena_b rc_osc_0.vr 0.746068f
C552 a_n10075_n19314# avss 0.466333f
C553 rstring_mux_0.vtrip_decoded_b_avdd[0] vin_vunder 0.269308f
C554 a_3748_n3212# rstring_mux_0.vtrip_decoded_avdd[2] 0.135857f
C555 rstring_mux_0.vtrip_decoded_avdd[6] avss 1.44633f
C556 a_n10463_9395# a_n9707_9395# 0.296258f
C557 rstring_mux_0.vtrip0 rstring_mux_0.vtrip2 0.847499f
C558 a_5346_n3990# avdd 0.607928f
C559 ibias_gen_0.vp1 avdd 6.59272f
C560 rstring_mux_0.vtrip_decoded_b_avdd[5] avss 0.363125f
C561 a_n8563_n19314# a_n7807_n19314# 0.296258f
C562 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_b_avdd[3] 0.571961f
C563 a_7033_n2212# avdd 0.142934f
C564 a_n26074_n2937# a_n25318_n2937# 0.296258f
C565 a_3911_n11914# a_4667_n11914# 0.296258f
C566 rstring_mux_0.otrip_decoded_avdd[6] dcomp3v3uv 0.148623f
C567 a_329_n1230# avdd 0.206171f
C568 rstring_mux_0.vtrip_decoded_b_avdd[6] avdd 0.904181f
C569 a_n15367_n19314# avss 0.466415f
C570 a_n6007_n2964# a_n5907_n2876# 0.40546f
C571 rstring_mux_0.otrip_decoded_b_avdd[1] avss 0.365652f
C572 a_10873_n3956# a_10514_n3890# 0.249269f
C573 a_329_n2964# dvdd 0.380879f
C574 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.vtrip4 0.192181f
C575 a_3748_n1478# rstring_mux_0.vtrip_decoded_avdd[3] 0.13699f
C576 a_n7429_n11914# vin_vunder 0.159467f
C577 rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.vtrip2 0.478934f
C578 comparator_0.vpp comparator_0.vnn 8.532559f
C579 rstring_mux_0.otrip_decoded_b_avdd[2] avdd 0.903648f
C580 sky130_fd_sc_hd__inv_4_1.Y dvdd 1.26215f
C581 ibias_gen_0.ena_b ibias_gen_0.isrc_sel_b 3.0701f
C582 comparator_0.vt comparator_0.vpp 2.58192f
C583 a_429_n2876# avdd 0.863791f
C584 comparator_1.n0 comparator_1.n1 0.927093f
C585 comparator_1.vnn comparator_1.vn 0.291139f
C586 comparator_1.vpp comparator_1.vm 0.633834f
C587 ibias_gen_0.ibias0 avdd 2.53198f
C588 rstring_mux_0.otrip_decoded_avdd[1] avdd 1.73956f
C589 a_n13855_n19314# a_n13099_n19314# 0.296258f
C590 a_5346_n2256# dvdd 0.104499f
C591 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[0] 0.260407f
C592 a_n8119_n2964# a_n7751_n3946# 0.138963f
C593 rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.vtrip4 0.533298f
C594 a_n6007_n1230# a_n5907_n1142# 0.40546f
C595 a_11121_n24601# a_11121_n25357# 0.296258f
C596 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y 0.392612f
C597 a_n12721_n11914# vin_vunder 0.159467f
C598 vl ibias_gen_0.isrc_sel 0.171708f
C599 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip_decoded_avdd[2] 1.78143f
C600 a_4553_n2964# vtrip_decoded[4] 0.2082f
C601 a_2809_n3946# dvdd 0.176016f
C602 rc_osc_0.in vin_vunder 0.174353f
C603 rstring_mux_0.vtrip4 avdd 0.416503f
C604 rstring_mux_0.otrip_decoded_avdd[0] dvdd 0.197825f
C605 a_n15479_n3901# ibg_200n 0.401026f
C606 a_10515_n1026# avdd 0.538412f
C607 dcomp3v3uv comparator_0.n0 0.388405f
C608 rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.vtrip6 0.489702f
C609 rstring_mux_0.vtrip_decoded_avdd[4] avss 1.50015f
C610 a_4921_n3946# avdd 0.143952f
C611 a_n8951_9395# avss 0.460284f
C612 a_3234_n3990# avdd 0.607928f
C613 rstring_mux_0.otrip_decoded_b_avdd[1] vin_brout 0.342078f
C614 rc_osc_0.m osc_ck 1.09227f
C615 comparator_1.vm avss 10.3557f
C616 a_n24562_n2937# avss 0.471605f
C617 a_n23428_n10337# a_n22672_n10337# 0.296258f
C618 dvdd outb_unbuf 0.331937f
C619 a_6557_n19314# a_7313_n19314# 0.296258f
C620 a_5423_n11914# avss 0.525451f
C621 a_9145_n2212# dvdd 0.169037f
C622 a_4553_n2964# a_4653_n2876# 0.40546f
C623 a_n8019_n2876# a_n7326_n3990# 0.264594f
C624 rstring_mux_0.vtrip_decoded_avdd[6] vin_vunder 0.880778f
C625 rstring_mux_0.vtrip0 rstring_mux_0.vtrip4 0.655814f
C626 dcomp3v3uv avdd 5.82321f
C627 a_n14243_9395# avss 0.460284f
C628 dvdd osc_ena 0.768954f
C629 rstring_mux_0.vtrip_decoded_b_avdd[5] vin_vunder 0.340862f
C630 a_n8185_n11914# a_n7429_n11914# 0.296258f
C631 a_n8119_n2964# avdd 0.194488f
C632 rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.otrip_decoded_b_avdd[2] 0.572197f
C633 a_131_n11914# avss 0.465554f
C634 ibias_gen_0.vp1 ibias_gen_0.isrc_sel 0.646099f
C635 a_1636_n1478# avdd 0.420074f
C636 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dcomp3v3uv 2.56892f
C637 a_n5907_n2876# a_n4700_n3212# 0.28899f
C638 a_n13109_1995# a_n12353_1995# 0.296258f
C639 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_avdd[2] 0.101824f
C640 comparator_0.ibias a_n27208_n10337# 0.311542f
C641 a_8069_n19314# avss 0.466333f
C642 a_n21916_n10337# avss 0.472978f
C643 a_3234_n2256# a_2809_n2212# 0.460766f
C644 a_8777_n1230# a_9145_n2212# 0.138963f
C645 sky130_fd_sc_hd__inv_4_4.Y dvdd 1.3053f
C646 rc_osc_0.in dvdd 5.53071f
C647 a_7972_n3212# rstring_mux_0.vtrip_decoded_avdd[6] 0.136133f
C648 a_1265_n19314# a_2021_n19314# 0.296258f
C649 a_n6673_n11914# avss 0.465068f
C650 a_3234_n2256# dvdd 0.104499f
C651 rstring_mux_0.otrip_decoded_b_avdd[6] avss 0.36281f
C652 a_4553_n1230# a_4653_n1142# 0.40546f
C653 a_n8019_n1142# a_n7326_n2256# 0.264594f
C654 comparator_0.vpp comparator_0.vn 0.332307f
C655 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip_decoded_avdd[2] 0.618116f
C656 a_n11597_1995# avss 0.460203f
C657 a_2441_n2964# avdd 0.207177f
C658 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip_decoded_b_avdd[3] 0.572316f
C659 comparator_1.n1 dcomp3v3 1.70353f
C660 comparator_1.vnn comparator_1.n0 0.42769f
C661 a_n27208_n10337# avss 0.761384f
C662 rstring_mux_0.otrip_decoded_b_avdd[7] avdd 0.903548f
C663 a_2777_n19314# avss 0.466333f
C664 comparator_1.vt comparator_1.vnn 4.17609f
C665 rstring_mux_0.vtrip_decoded_avdd[7] avdd 1.81913f
C666 a_n13477_n11914# a_n12721_n11914# 0.296258f
C667 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[6] 0.211299f
C668 a_10874_n1026# dvdd 0.443515f
C669 comparator_0.ibias comparator_0.vnn 0.116472f
C670 a_n11965_n11914# avss 0.465068f
C671 rstring_mux_0.vtrip_decoded_avdd[2] avss 1.41004f
C672 a_n5907_n1142# a_n4700_n1478# 0.28899f
C673 a_n8119_n1230# dvdd 0.387414f
C674 rc_osc_0.in a_n10279_n24979# 0.770709f
C675 a_1122_n3990# avdd 0.607928f
C676 a_2441_n1230# vtrip_decoded[3] 0.2082f
C677 rstring_mux_0.vtrip6 avdd 0.949337f
C678 rstring_mux_0.vtrip_decoded_avdd[6] dvdd 0.309916f
C679 a_7458_n2256# avdd 0.607928f
C680 vl rstring_mux_0.otrip_decoded_avdd[1] 0.145098f
C681 comparator_1.vn avdd 0.751908f
C682 a_7972_n1478# rstring_mux_0.vtrip_decoded_avdd[7] 0.13699f
C683 a_n4027_n19314# avss 0.466333f
C684 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.vtrip2 0.190544f
C685 rstring_mux_0.otrip_decoded_avdd[2] dcomp3v3uv 0.375655f
C686 a_n8019_n1142# avdd 0.864468f
C687 a_7033_n3946# avdd 0.143952f
C688 rstring_mux_0.vtrip_decoded_avdd[4] vin_vunder 0.875594f
C689 a_n5539_n19314# a_n4783_n19314# 0.296258f
C690 comparator_0.vnn avss 3.54397f
C691 a_n23050_n2937# a_n22294_n2937# 0.296258f
C692 comparator_1.n1 avss 2.99005f
C693 a_n990_n2256# a_n1415_n2212# 0.460766f
C694 a_6935_n11914# a_7691_n11914# 0.296258f
C695 comparator_0.vt avss 29.296902f
C696 rstring_mux_0.otrip_decoded_b_avdd[6] vin_brout 0.340862f
C697 a_2441_n1230# a_2809_n2212# 0.138963f
C698 rstring_mux_0.vtrip0 a_n4405_n11914# 0.137908f
C699 a_10873_n2760# a_10873_n3956# 0.136815f
C700 a_n9319_n19314# avss 0.466333f
C701 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_b_avdd[6] 0.155152f
C702 a_4653_n2876# a_5860_n3212# 0.28899f
C703 a_2441_n1230# dvdd 0.379209f
C704 rstring_mux_0.vtrip2 rstring_mux_0.vtrip4 0.994518f
C705 a_n6812_n3212# avdd 0.421965f
C706 comparator_0.ena a_n27208_n10337# 0.294281f
C707 a_131_n11914# vin_vunder 0.329686f
C708 a_2541_n1142# avdd 0.863296f
C709 a_1122_n2256# dvdd 0.104499f
C710 rc_osc_0.vr osc_ck 0.639788f
C711 a_n14611_n19314# avss 0.466333f
C712 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip_decoded_avdd[0] 1.27051f
C713 a_n12731_9395# a_n11975_9395# 0.296258f
C714 a_n10831_n19314# a_n10075_n19314# 0.296258f
C715 rstring_mux_0.vtrip_decoded_avdd[5] avdd 2.25645f
C716 a_1643_n11914# a_2399_n11914# 0.296258f
C717 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[4] 0.158489f
C718 a_4653_n1142# a_5860_n1478# 0.28899f
C719 a_n6673_n11914# vin_vunder 0.159467f
C720 comparator_0.ena_b comparator_0.vn 1.12681f
C721 comparator_0.vnn comparator_0.vm 0.573444f
C722 comparator_0.vpp comparator_0.n0 0.356806f
C723 a_n3795_n2876# a_n3102_n3990# 0.264594f
C724 rstring_mux_0.vtrip_decoded_avdd[0] avss 1.37856f
C725 a_n990_n3990# avdd 0.607928f
C726 ibias_gen_0.ena_b a_n15529_n2223# 0.244191f
C727 rstring_mux_0.vtrip_decoded_b_avdd[3] avss 0.362811f
C728 comparator_0.ena comparator_0.vnn 0.503016f
C729 a_3748_n3212# avdd 0.421965f
C730 rstring_mux_0.vtrip_decoded_avdd[4] dvdd 0.669746f
C731 rstring_mux_0.vtrip_decoded_avdd[2] rstring_mux_0.vtrip_decoded_b_avdd[2] 0.5727f
C732 a_n5214_n2256# a_n5639_n2212# 0.460766f
C733 a_5346_n3990# a_4921_n3946# 0.460766f
C734 comparator_1.vpp comparator_1.vnn 8.65712f
C735 sky130_fd_sc_hd__inv_4_3.Y dvdd 1.31104f
C736 a_6665_n2964# vtrip_decoded[6] 0.207265f
C737 a_9570_n2256# dvdd 0.103732f
C738 a_n6007_n2964# a_n5639_n3946# 0.138963f
C739 rstring_mux_0.vtrip_decoded_b_avdd[4] avdd 0.903548f
C740 comparator_0.ibias comparator_0.vn 0.423513f
C741 a_n11965_n11914# vin_vunder 0.159467f
C742 rstring_mux_0.vtrip_decoded_avdd[2] vin_vunder 0.884578f
C743 a_9145_n3946# dvdd 0.17571f
C744 comparator_0.vpp avdd 37.2833f
C745 comparator_1.n0 avdd 0.973197f
C746 a_10874_n2222# avdd 0.258197f
C747 comparator_1.vt avdd 0.141755p
C748 a_n3795_n1142# a_n3102_n2256# 0.264594f
C749 ibias_gen_0.vp1 dcomp3v3uv 0.195418f
C750 a_n6007_n1230# avdd 0.206171f
C751 a_n16123_n19314# a_n15367_n19314# 0.296258f
C752 rstring_mux_0.otrip_decoded_b_avdd[0] avdd 0.870606f
C753 a_n8195_9395# avss 0.721623f
C754 a_n5161_n11914# a_n4405_n11914# 0.296258f
C755 a_11121_n22333# a_11121_n23089# 0.296258f
C756 comparator_0.vn avss 8.8444f
C757 comparator_0.vnn vin_vunder 3.10064f
C758 a_n23806_n2937# avss 0.474081f
C759 comparator_1.vnn avss 3.08013f
C760 a_6179_n11914# avss 0.525451f
C761 comparator_0.vt vin_vunder 25.477098f
C762 a_n6007_n2964# dvdd 0.380879f
C763 a_6765_n2876# a_7458_n3990# 0.264594f
C764 a_n990_n2256# dvdd 0.104499f
C765 rstring_mux_0.vtrip_decoded_avdd[0] vin_brout 0.252789f
C766 a_n10085_1995# a_n9329_1995# 0.296258f
C767 rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.otrip_decoded_b_avdd[5] 0.155092f
C768 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.vtrip_decoded_avdd[0] 0.34246f
C769 a_n13487_9395# avss 0.460203f
C770 vl a_n14621_1995# 0.308117f
C771 a_n5907_n2876# avdd 0.863791f
C772 a_n25696_n10337# a_n24940_n10337# 0.296258f
C773 rstring_mux_0.vtrip_decoded_avdd[3] avdd 1.87754f
C774 a_1122_n3990# a_697_n3946# 0.460766f
C775 a_887_n11914# avss 0.465525f
C776 a_4289_n19314# a_5045_n19314# 0.296258f
C777 a_4553_n1230# avdd 0.206171f
C778 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.vtrip0 0.191117f
C779 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[2] 0.13771f
C780 sky130_fd_sc_hd__inv_4_4.Y outb_unbuf 0.396003f
C781 rstring_mux_0.otrip_decoded_avdd[6] avss 1.36421f
C782 a_n3895_n2964# a_n3795_n2876# 0.40546f
C783 a_n3102_n3990# avdd 0.607928f
C784 a_8825_n19314# avss 0.466415f
C785 a_n21160_n10337# avss 0.476371f
C786 a_10873_n2760# dvdd 0.443538f
C787 rstring_mux_0.vtrip_decoded_avdd[2] dvdd 0.279976f
C788 a_n10453_n11914# a_n9697_n11914# 0.296258f
C789 a_4553_n2964# dvdd 0.380879f
C790 a_n5917_n11914# avss 0.465068f
C791 rstring_mux_0.vtrip_decoded_avdd[7] rstring_mux_0.vtrip_decoded_b_avdd[6] 0.155139f
C792 rc_osc_0.in osc_ena 0.161388f
C793 schmitt_trigger_0.in comparator_0.vnn 0.268371f
C794 comparator_0.vn comparator_0.vm 4.66142f
C795 rstring_mux_0.vtrip_decoded_avdd[0] vin_vunder 0.599238f
C796 a_7458_n3990# avdd 0.607928f
C797 a_n10841_1995# avss 0.460203f
C798 comparator_1.vnn vin_brout 2.4293f
C799 comparator_0.ena comparator_0.vn 0.139186f
C800 rstring_mux_0.vtrip_decoded_b_avdd[3] vin_vunder 0.340862f
C801 a_4653_n2876# avdd 0.863791f
C802 a_7458_n2256# a_7033_n2212# 0.460766f
C803 a_n8119_n2964# otrip_decoded[0] 0.207169f
C804 a_3533_n19314# avss 0.466333f
C805 a_n26452_n10337# avss 0.47306f
C806 a_10514_n2760# a_10514_n3890# 0.170258f
C807 comparator_1.vnn comparator_0.ena 0.731104f
C808 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip6 0.190544f
C809 rstring_mux_0.ena_b avss 1.61845f
C810 a_4553_n1230# vtrip_decoded[5] 0.2082f
C811 a_n7751_n2212# dvdd 0.169579f
C812 a_n3895_n1230# a_n3795_n1142# 0.40546f
C813 a_n11209_n11914# avss 0.465068f
C814 a_n9319_n19314# dvdd 0.407976f
C815 avdd itest 0.241333f
C816 comparator_0.ena_b avdd 1.01938f
C817 dcomp3v3 avdd 6.72634f
C818 a_n5639_n2212# avdd 0.142934f
C819 comparator_1.vpp avdd 37.1895f
C820 a_n3102_n3990# a_n3527_n3946# 0.460766f
C821 a_n4700_n1478# avdd 0.420074f
C822 rstring_mux_0.otrip_decoded_b_avdd[4] avss 0.36282f
C823 rstring_mux_0.otrip_decoded_avdd[6] vin_brout 0.875633f
C824 a_429_n2876# a_1122_n3990# 0.264594f
C825 a_n3102_n2256# dvdd 0.104499f
C826 a_n15745_n11914# a_n14989_n11914# 0.296258f
C827 comparator_0.n0 avss 4.20459f
C828 a_n10279_n22711# a_n10279_n23467# 0.296258f
C829 comparator_0.ibias avdd 7.48627f
C830 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_avdd[6] 1.12965f
C831 vl a_10874_n2222# 0.153476f
C832 rstring_mux_0.otrip_decoded_b_avdd[5] avdd 0.903548f
C833 ibias_gen_0.ibias0 comparator_1.vn 0.59661f
C834 rstring_mux_0.vtrip0 a_n3649_n11914# 0.411488f
C835 a_4553_n1230# a_4921_n2212# 0.138963f
C836 rc_osc_0.m dvdd 2.38628f
C837 rstring_mux_0.vtrip_decoded_avdd[1] avdd 1.96911f
C838 schmitt_trigger_0.in rstring_mux_0.vtrip_decoded_avdd[0] 0.128751f
C839 a_n8563_n19314# avss 0.466333f
C840 a_n9707_9395# a_n8951_9395# 0.296258f
C841 a_6665_n2964# a_6765_n2876# 0.40546f
C842 rstring_mux_0.otrip_decoded_avdd[4] avss 1.34995f
C843 rstring_mux_0.vtrip4 rstring_mux_0.vtrip6 0.859994f
C844 a_n5214_n3990# avdd 0.607928f
C845 a_n7807_n19314# a_n7051_n19314# 0.296258f
C846 a_n3895_n2964# avdd 0.207177f
C847 avdd avss 2.43878p
C848 rstring_mux_0.vtrip_decoded_avdd[0] dvdd 0.275187f
C849 a_n25318_n2937# a_n24562_n2937# 0.296258f
C850 a_4667_n11914# a_5423_n11914# 0.296258f
C851 a_429_n1142# a_1122_n2256# 0.264594f
C852 a_5860_n1478# avdd 0.420074f
C853 comparator_0.ena rstring_mux_0.ena_b 0.179228f
C854 a_n13855_n19314# avss 0.466333f
C855 a_n3795_n2876# a_n2588_n3212# 0.28899f
C856 a_9570_n3990# dvdd 0.103731f
C857 a_n14999_9395# avss 0.721623f
C858 avss ibg_200n 0.598217f
C859 rstring_mux_0.otrip_decoded_b_avdd[4] vin_brout 0.340862f
C860 a_n7326_n3990# a_n7751_n3946# 0.460766f
C861 a_6665_n1230# a_6765_n1142# 0.40546f
C862 a_n5917_n11914# vin_vunder 0.159467f
C863 rstring_mux_0.vtrip_decoded_avdd[6] rstring_mux_0.vtrip_decoded_b_avdd[5] 0.155037f
C864 comparator_0.vm comparator_0.n0 2.61558f
C865 a_10873_n3956# avdd 0.258162f
C866 a_8777_n2964# ena 0.2082f
C867 rstring_mux_0.vtrip0 avss 2.36542f
C868 a_9570_n2256# a_9145_n2212# 0.460766f
C869 a_6665_n2964# avdd 0.207177f
C870 a_n3527_n2212# dvdd 0.169343f
C871 a_n13099_n19314# a_n12343_n19314# 0.296258f
C872 a_n5214_n2256# dvdd 0.105303f
C873 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X a_10873_n3956# 0.142786f
C874 a_n3895_n2964# a_n3527_n3946# 0.138963f
C875 rstring_mux_0.otrip_decoded_avdd[4] vin_brout 0.879587f
C876 a_n3795_n1142# a_n2588_n1478# 0.28899f
C877 a_n11209_n11914# vin_vunder 0.159467f
C878 a_n3895_n1230# dvdd 0.38629f
C879 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_avdd[6] 0.340239f
C880 comparator_0.vm avdd 0.390636f
C881 avdd vin_brout 6.34191f
C882 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip_decoded_b_avdd[1] 0.572131f
C883 a_n1415_n2212# avdd 0.142934f
C884 rstring_mux_0.ena_b rstring_mux_0.vtop 2.52783f
C885 comparator_0.ena avdd 17.5497f
C886 sky130_fd_sc_hd__inv_4_0.Y dvdd 1.35239f
C887 rstring_mux_0.otrip_decoded_avdd[7] avdd 1.82047f
C888 a_n3795_n1142# avdd 0.863296f
C889 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[6] 0.105908f
C890 dcomp3v3 ibias_gen_0.isrc_sel 10.963901f
C891 rstring_mux_0.otrip_decoded_avdd[2] avss 1.41238f
C892 comparator_0.n0 vin_vunder 0.103885f
C893 rstring_mux_0.vtrip_decoded_b_avdd[1] avss 0.362828f
C894 a_n7326_n3990# avdd 0.607831f
C895 a_6935_n11914# avss 0.525451f
C896 a_n22672_n10337# a_n21916_n10337# 0.296258f
C897 a_n23050_n2937# avss 0.474704f
C898 dcomp3v3 vl 10.054f
C899 rstring_mux_0.otrip_decoded_avdd[6] dvdd 0.257138f
C900 a_7313_n19314# a_8069_n19314# 0.296258f
C901 ibias_gen_0.ibias0 comparator_1.n0 0.172673f
C902 dvdd dcomp 1.54533f
C903 comparator_1.vt ibias_gen_0.ibias0 0.504592f
C904 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip4 0.190544f
C905 comparator_0.ena ibg_200n 0.218863f
C906 a_8877_n2876# a_9570_n3990# 0.264594f
C907 a_6665_n1230# dvdd 0.379209f
C908 a_n2588_n3212# rstring_mux_0.otrip_decoded_avdd[4] 0.136088f
C909 a_6765_n2876# a_7972_n3212# 0.28899f
C910 rstring_mux_0.vtrip0 vin_brout 2.24047f
C911 rstring_mux_0.vtrip_decoded_b_avdd[2] avdd 0.903548f
C912 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_b_avdd[0] 0.176375f
C913 vl comparator_0.ibias 0.261037f
C914 a_n12731_9395# avss 0.460203f
C915 a_n7429_n11914# a_n6673_n11914# 0.296258f
C916 a_n2588_n3212# avdd 0.421965f
C917 a_10515_n1026# a_10874_n2222# 0.166612f
C918 comparator_0.vnn vbg_1v2 0.779817f
C919 a_1643_n11914# avss 0.465635f
C920 a_10514_n2760# a_10873_n2760# 0.249533f
C921 avdd vin_vunder 5.50314f
C922 comparator_0.vt vbg_1v2 24.362598f
C923 a_6765_n1142# avdd 0.863296f
C924 a_4653_n2876# a_5346_n3990# 0.264594f
C925 ibias_gen_0.isrc_sel avss 3.29158f
C926 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_b_avdd[4] 0.155007f
C927 a_n12353_1995# a_n11597_1995# 0.296258f
C928 rc_osc_0.vr dvdd 1.51499f
C929 a_n20404_n10337# avss 0.769579f
C930 a_n7751_n3946# dvdd 0.176029f
C931 a_9581_n19314# avss 0.730849f
C932 vl avss 1.65817f
C933 rstring_mux_0.vtop avdd 10.640901f
C934 rstring_mux_0.vtrip6 a_n247_n19314# 0.298448f
C935 a_n5161_n11914# avss 0.475109f
C936 a_n2588_n1478# rstring_mux_0.otrip_decoded_avdd[5] 0.13699f
C937 a_2021_n19314# a_2777_n19314# 0.296258f
C938 a_6765_n1142# a_7972_n1478# 0.28899f
C939 a_n7326_n2256# dvdd 0.104499f
C940 rstring_mux_0.otrip_decoded_avdd[2] vin_brout 0.880848f
C941 comparator_0.n0 comparator_0.n1 0.927063f
C942 a_n6007_n2964# otrip_decoded[2] 0.2082f
C943 dcomp3v3 ibias_gen_0.vp1 0.543408f
C944 a_n5639_n3946# avdd 0.145138f
C945 a_n10085_1995# avss 0.460203f
C946 rstring_mux_0.vtrip2 avss 2.19733f
C947 a_6665_n1230# vtrip_decoded[7] 0.2082f
C948 rstring_mux_0.vtrip0 vin_vunder 2.24424f
C949 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_avdd[4] 1.15427f
C950 a_7972_n3212# avdd 0.421965f
C951 a_n25696_n10337# avss 0.472978f
C952 a_4289_n19314# avss 0.466333f
C953 sky130_fd_sc_hd__inv_4_0.Y brout_filt 1.46398f
C954 a_4653_n1142# a_5346_n2256# 0.264594f
C955 a_697_n2212# dvdd 0.169343f
C956 rstring_mux_0.otrip_decoded_avdd[5] avdd 1.82417f
C957 a_n12721_n11914# a_n11965_n11914# 0.296258f
C958 ibias_gen_0.vp1 comparator_0.ibias 0.404784f
C959 a_n10453_n11914# avss 0.465068f
C960 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[4] 0.101976f
C961 schmitt_trigger_0.in avdd 3.79238f
C962 comparator_0.n1 avdd 2.68846f
C963 rstring_mux_0.otrip_decoded_avdd[4] dvdd 0.266092f
C964 rstring_mux_0.vtrip_decoded_avdd[0] rstring_mux_0.vtrip_decoded_b_avdd[0] 0.574058f
C965 a_2809_n2212# avdd 0.142934f
C966 a_n1783_n1230# avdd 0.206171f
C967 avdd dvdd 42.420998f
C968 ibias_gen_0.vp1 avss 2.02475f
C969 a_n15745_n11914# avss 0.465267f
C970 a_n4783_n19314# a_n4027_n19314# 0.296258f
C971 comparator_0.ena ibias_gen_0.isrc_sel 1.49913f
C972 rstring_mux_0.vtrip_decoded_b_avdd[1] vin_vunder 0.340862f
C973 a_n22294_n2937# a_n21538_n2937# 0.296258f
C974 a_7691_n11914# a_8447_n11914# 0.296258f
C975 comparator_0.vt rc_osc_0.in 0.164658f
C976 comparator_1.vpp ibias_gen_0.ibias0 1.31426f
C977 a_n1783_n2964# dvdd 0.380879f
C978 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd 1.32384f
C979 rstring_mux_0.vtrip_decoded_b_avdd[6] avss 0.363573f
C980 a_n7807_n19314# avss 0.466333f
C981 rc_osc_0.m osc_ena 0.252626f
C982 rstring_mux_0.vtrip2 vin_brout 2.09579f
C983 ibias_gen_0.ena_b avdd 2.96986f
C984 dcomp3v3 a_10515_n1026# 0.207687f
C985 a_n1683_n2876# avdd 0.863791f
C986 rstring_mux_0.vtrip_decoded_b_avdd[7] avdd 0.839308f
C987 comparator_0.vn vbg_1v2 0.728008f
C988 comparator_1.vn comparator_1.n0 1.97873f
C989 comparator_1.vt comparator_1.vn 0.203925f
C990 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X sky130_fd_sc_hd__inv_4_1.A 0.431807f
C991 a_8777_n1230# avdd 0.206179f
C992 comparator_1.vnn vbg_1v2 1.97725f
C993 a_n8119_n1230# a_n7751_n2212# 0.138963f
C994 osc_ck dvss 3.25723f
C995 osc_ena dvss 2.21578f
C996 vin_vunder dvss 42.69882f
C997 ena dvss 0.377679f
C998 vtrip_decoded[6] dvss 0.373773f
C999 vtrip_decoded[4] dvss 0.377387f
C1000 vtrip_decoded[2] dvss 0.37758f
C1001 vtrip_decoded[0] dvss 0.37744f
C1002 otrip_decoded[6] dvss 0.378276f
C1003 otrip_decoded[4] dvss 0.384187f
C1004 otrip_decoded[2] dvss 0.382228f
C1005 otrip_decoded[0] dvss 0.403289f
C1006 isrc_sel dvss 0.383453f
C1007 vtrip_decoded[7] dvss 0.375086f
C1008 vtrip_decoded[5] dvss 0.375086f
C1009 vtrip_decoded[3] dvss 0.375086f
C1010 vtrip_decoded[1] dvss 0.375086f
C1011 otrip_decoded[7] dvss 0.375086f
C1012 otrip_decoded[5] dvss 0.373107f
C1013 otrip_decoded[3] dvss 0.372167f
C1014 otrip_decoded[1] dvss 0.397873f
C1015 vunder dvss 1.25924f
C1016 brout_filt dvss 1.31887f
C1017 dcomp dvss 1.25747f
C1018 outb dvss 1.26961f
C1019 outb_unbuf dvss 0.626298f
C1020 ibg_200n dvss 0.16009f
C1021 itest dvss 0.296385f
C1022 vbg_1v2 dvss 47.65465f
C1023 vin_brout dvss 24.391699f
C1024 dvdd dvss 1.0343p
C1025 avss dvss 0.211383p
C1026 avdd dvss 3.602057p
C1027 a_11121_n25357# dvss 1.41754f
C1028 a_n10279_n24979# dvss 1.13069f
C1029 a_11121_n24601# dvss 1.13097f
C1030 a_n10279_n24223# dvss 1.13821f
C1031 a_11121_n23845# dvss 1.13089f
C1032 a_n10279_n23467# dvss 1.31493f
C1033 a_11121_n23089# dvss 1.13097f
C1034 a_n10279_n22711# dvss 1.20647f
C1035 a_11121_n22333# dvss 1.398f
C1036 rc_osc_0.vr dvss 4.10332f
C1037 rc_osc_0.m dvss 3.35349f
C1038 rc_osc_0.in dvss 0.439754p
C1039 rc_osc_0.ena_b dvss 1.39535f
C1040 a_9581_n19314# dvss 0.612822f
C1041 a_9203_n11914# dvss 0.659772f
C1042 a_8825_n19314# dvss 0.61321f
C1043 a_8447_n11914# dvss 0.659772f
C1044 a_8069_n19314# dvss 0.61321f
C1045 a_7691_n11914# dvss 0.659772f
C1046 a_7313_n19314# dvss 0.61321f
C1047 a_6935_n11914# dvss 0.659772f
C1048 a_6557_n19314# dvss 0.61321f
C1049 a_6179_n11914# dvss 0.659772f
C1050 a_5801_n19314# dvss 0.61321f
C1051 a_5423_n11914# dvss 0.659772f
C1052 a_5045_n19314# dvss 0.618291f
C1053 a_4667_n11914# dvss 0.659772f
C1054 a_4289_n19314# dvss 0.61321f
C1055 a_3911_n11914# dvss 0.647659f
C1056 a_3533_n19314# dvss 0.61321f
C1057 a_3155_n11914# dvss 0.653638f
C1058 a_2777_n19314# dvss 0.61321f
C1059 a_2399_n11914# dvss 0.656775f
C1060 a_2021_n19314# dvss 0.61321f
C1061 a_1643_n11914# dvss 0.656775f
C1062 a_1265_n19314# dvss 0.61321f
C1063 a_887_n11914# dvss 0.656775f
C1064 a_509_n19314# dvss 0.61321f
C1065 a_131_n11914# dvss 0.642157f
C1066 a_n247_n19314# dvss 0.61321f
C1067 a_n3649_n11914# dvss 0.635008f
C1068 a_n4027_n19314# dvss 0.61321f
C1069 a_n4405_n11914# dvss 0.640419f
C1070 a_n4783_n19314# dvss 0.61321f
C1071 a_n5161_n11914# dvss 0.643911f
C1072 a_n5539_n19314# dvss 0.61321f
C1073 a_n5917_n11914# dvss 0.643911f
C1074 a_n6295_n19314# dvss 0.61321f
C1075 a_n6673_n11914# dvss 0.643911f
C1076 a_n7051_n19314# dvss 0.61321f
C1077 a_n7429_n11914# dvss 0.645008f
C1078 a_n7807_n19314# dvss 0.621617f
C1079 a_n8185_n11914# dvss 0.651324f
C1080 a_n8563_n19314# dvss 0.644889f
C1081 a_n8941_n11914# dvss 1.04349f
C1082 a_n9319_n19314# dvss 0.978123f
C1083 a_n9697_n11914# dvss 0.626761f
C1084 a_n10075_n19314# dvss 0.61321f
C1085 a_n10453_n11914# dvss 0.643911f
C1086 a_n10831_n19314# dvss 0.61321f
C1087 a_n11209_n11914# dvss 0.643911f
C1088 a_n11587_n19314# dvss 0.61321f
C1089 a_n11965_n11914# dvss 0.643911f
C1090 a_n12343_n19314# dvss 0.61321f
C1091 a_n12721_n11914# dvss 0.643911f
C1092 a_n13099_n19314# dvss 0.61321f
C1093 a_n13477_n11914# dvss 0.643911f
C1094 a_n13855_n19314# dvss 0.612139f
C1095 a_n14233_n11914# dvss 0.643911f
C1096 a_n14611_n19314# dvss 0.615216f
C1097 a_n14989_n11914# dvss 0.643911f
C1098 a_n15367_n19314# dvss 0.61321f
C1099 a_n15745_n11914# dvss 0.628722f
C1100 a_n16123_n19314# dvss 0.612803f
C1101 comparator_0.n1 dvss 1.57269f
C1102 comparator_0.n0 dvss 0.809097f
C1103 comparator_0.vm dvss 4.68965f
C1104 comparator_0.vn dvss 5.29407f
C1105 comparator_0.ena_b dvss 0.795107f
C1106 comparator_0.vnn dvss 44.4198f
C1107 comparator_0.vpp dvss 38.2285f
C1108 rstring_mux_0.vtrip6 dvss 6.108224f
C1109 rstring_mux_0.vtrip4 dvss 5.681643f
C1110 rstring_mux_0.vtrip2 dvss 5.372343f
C1111 rstring_mux_0.vtrip0 dvss 7.09113f
C1112 rstring_mux_0.vtop dvss 16.18401f
C1113 rstring_mux_0.ena_b dvss 2.14258f
C1114 rstring_mux_0.vtrip_decoded_b_avdd[7] dvss 0.214336f
C1115 rstring_mux_0.vtrip_decoded_b_avdd[6] dvss 0.191802f
C1116 rstring_mux_0.vtrip_decoded_b_avdd[5] dvss 0.191802f
C1117 rstring_mux_0.vtrip_decoded_b_avdd[4] dvss 0.191802f
C1118 rstring_mux_0.vtrip_decoded_b_avdd[3] dvss 0.191802f
C1119 rstring_mux_0.vtrip_decoded_b_avdd[2] dvss 0.191802f
C1120 rstring_mux_0.vtrip_decoded_b_avdd[1] dvss 0.191801f
C1121 rstring_mux_0.vtrip_decoded_b_avdd[0] dvss 0.193218f
C1122 rstring_mux_0.otrip_decoded_b_avdd[7] dvss 0.191802f
C1123 rstring_mux_0.otrip_decoded_b_avdd[6] dvss 0.191802f
C1124 rstring_mux_0.otrip_decoded_b_avdd[5] dvss 0.191802f
C1125 rstring_mux_0.otrip_decoded_b_avdd[4] dvss 0.191802f
C1126 rstring_mux_0.otrip_decoded_b_avdd[3] dvss 0.181122f
C1127 rstring_mux_0.otrip_decoded_b_avdd[2] dvss 0.191802f
C1128 rstring_mux_0.otrip_decoded_b_avdd[1] dvss 0.191802f
C1129 rstring_mux_0.otrip_decoded_b_avdd[0] dvss 0.195093f
C1130 a_9145_n3946# dvss 1.70782f
C1131 a_7033_n3946# dvss 1.70837f
C1132 a_10514_n3890# dvss 0.90142f
C1133 a_4921_n3946# dvss 1.70837f
C1134 a_2809_n3946# dvss 1.70837f
C1135 a_697_n3946# dvss 1.70837f
C1136 a_n1415_n3946# dvss 1.70837f
C1137 a_n3527_n3946# dvss 1.70837f
C1138 a_n5639_n3946# dvss 1.70837f
C1139 a_n7751_n3946# dvss 1.70982f
C1140 a_10873_n3956# dvss 1.0124f
C1141 a_9570_n3990# dvss 0.849936f
C1142 a_7458_n3990# dvss 0.867563f
C1143 a_10873_n2760# dvss 0.860482f
C1144 dcomp3v3uv dvss 7.377871f
C1145 a_10514_n2760# dvss 1.27441f
C1146 a_5346_n3990# dvss 0.867571f
C1147 rstring_mux_0.vtrip_decoded_avdd[6] dvss 1.45409f
C1148 a_3234_n3990# dvss 0.867563f
C1149 rstring_mux_0.vtrip_decoded_avdd[4] dvss 1.43527f
C1150 a_1122_n3990# dvss 0.867563f
C1151 rstring_mux_0.vtrip_decoded_avdd[2] dvss 1.70338f
C1152 a_n990_n3990# dvss 0.867563f
C1153 rstring_mux_0.vtrip_decoded_avdd[0] dvss 1.48566f
C1154 a_n3102_n3990# dvss 0.867563f
C1155 rstring_mux_0.otrip_decoded_avdd[6] dvss 1.25006f
C1156 a_n5214_n3990# dvss 0.867563f
C1157 rstring_mux_0.otrip_decoded_avdd[4] dvss 1.06381f
C1158 a_n7326_n3990# dvss 0.867659f
C1159 rstring_mux_0.otrip_decoded_avdd[2] dvss 1.43078f
C1160 rstring_mux_0.otrip_decoded_avdd[0] dvss 1.07955f
C1161 a_10084_n3212# dvss 0.492184f
C1162 a_8877_n2876# dvss 1.52129f
C1163 a_8777_n2964# dvss 1.97869f
C1164 a_7972_n3212# dvss 0.503164f
C1165 a_6765_n2876# dvss 1.52226f
C1166 a_6665_n2964# dvss 1.97975f
C1167 a_5860_n3212# dvss 0.503164f
C1168 a_4653_n2876# dvss 1.52226f
C1169 a_4553_n2964# dvss 1.97975f
C1170 a_3748_n3212# dvss 0.503164f
C1171 a_2541_n2876# dvss 1.52226f
C1172 a_2441_n2964# dvss 1.97975f
C1173 a_1636_n3212# dvss 0.503164f
C1174 a_429_n2876# dvss 1.52226f
C1175 a_329_n2964# dvss 1.97975f
C1176 a_n476_n3212# dvss 0.503164f
C1177 a_n1683_n2876# dvss 1.52226f
C1178 a_n1783_n2964# dvss 1.97975f
C1179 a_n2588_n3212# dvss 0.503164f
C1180 a_n3795_n2876# dvss 1.52226f
C1181 a_n3895_n2964# dvss 1.97975f
C1182 a_n4700_n3212# dvss 0.503164f
C1183 a_n5907_n2876# dvss 1.52226f
C1184 a_n6007_n2964# dvss 1.97975f
C1185 a_n6812_n3212# dvss 0.503164f
C1186 a_n8019_n2876# dvss 1.53095f
C1187 a_n8119_n2964# dvss 2.03637f
C1188 a_9145_n2212# dvss 1.69093f
C1189 a_7033_n2212# dvss 1.69148f
C1190 a_10515_n2156# dvss 0.891723f
C1191 a_4921_n2212# dvss 1.69148f
C1192 a_2809_n2212# dvss 1.69148f
C1193 a_697_n2212# dvss 1.69148f
C1194 a_n1415_n2212# dvss 1.69148f
C1195 a_n3527_n2212# dvss 1.69148f
C1196 a_n5639_n2212# dvss 1.69215f
C1197 a_n7751_n2212# dvss 1.69294f
C1198 a_10874_n2222# dvss 1.00525f
C1199 a_9570_n2256# dvss 0.84998f
C1200 a_7458_n2256# dvss 0.867563f
C1201 a_10874_n1026# dvss 0.862185f
C1202 a_10515_n1026# dvss 1.27471f
C1203 a_5346_n2256# dvss 0.867563f
C1204 rstring_mux_0.vtrip_decoded_avdd[7] dvss 2.19103f
C1205 a_3234_n2256# dvss 0.867563f
C1206 rstring_mux_0.vtrip_decoded_avdd[5] dvss 1.9559f
C1207 a_1122_n2256# dvss 0.867563f
C1208 rstring_mux_0.vtrip_decoded_avdd[3] dvss 2.02174f
C1209 a_n990_n2256# dvss 0.867563f
C1210 rstring_mux_0.vtrip_decoded_avdd[1] dvss 2.11486f
C1211 a_n3102_n2256# dvss 0.867563f
C1212 rstring_mux_0.otrip_decoded_avdd[7] dvss 1.87654f
C1213 a_n5214_n2256# dvss 0.867974f
C1214 rstring_mux_0.otrip_decoded_avdd[5] dvss 1.92238f
C1215 a_n7326_n2256# dvss 0.867659f
C1216 rstring_mux_0.otrip_decoded_avdd[3] dvss 1.59657f
C1217 rstring_mux_0.otrip_decoded_avdd[1] dvss 1.75829f
C1218 a_10084_n1478# dvss 0.490437f
C1219 a_8877_n1142# dvss 1.52856f
C1220 a_8777_n1230# dvss 1.97228f
C1221 a_7972_n1478# dvss 0.501383f
C1222 a_6765_n1142# dvss 1.52953f
C1223 a_6665_n1230# dvss 1.97335f
C1224 a_5860_n1478# dvss 0.501383f
C1225 a_4653_n1142# dvss 1.52953f
C1226 a_4553_n1230# dvss 1.97335f
C1227 a_3748_n1478# dvss 0.501383f
C1228 a_2541_n1142# dvss 1.52953f
C1229 a_2441_n1230# dvss 1.97335f
C1230 a_1636_n1478# dvss 0.501383f
C1231 a_429_n1142# dvss 1.52953f
C1232 a_329_n1230# dvss 1.97335f
C1233 a_n476_n1478# dvss 0.501383f
C1234 a_n1683_n1142# dvss 1.52953f
C1235 a_n1783_n1230# dvss 1.96643f
C1236 a_n2588_n1478# dvss 0.500163f
C1237 a_n3795_n1142# dvss 1.52683f
C1238 a_n3895_n1230# dvss 1.96734f
C1239 a_n4700_n1478# dvss 0.512534f
C1240 a_n5907_n1142# dvss 1.53695f
C1241 a_n6007_n1230# dvss 1.97338f
C1242 a_n6812_n1478# dvss 0.501043f
C1243 a_n8019_n1142# dvss 1.53771f
C1244 a_n8119_n1230# dvss 2.02842f
C1245 sky130_fd_sc_hd__inv_4_1.Y dvss 2.05205f
C1246 sky130_fd_sc_hd__inv_4_1.A dvss 0.780068f
C1247 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss 4.01021f
C1248 sky130_fd_sc_hd__inv_4_0.Y dvss 1.95792f
C1249 schmitt_trigger_0.m dvss 2.365713f
C1250 sky130_fd_sc_hd__inv_4_3.Y dvss 1.98879f
C1251 sky130_fd_sc_hd__inv_4_4.Y dvss 2.01806f
C1252 a_n20404_n10337# dvss 0.639031f
C1253 a_n20782_n2937# dvss 0.502711f
C1254 a_n21160_n10337# dvss 0.639742f
C1255 a_n21538_n2937# dvss 0.502711f
C1256 a_n21916_n10337# dvss 0.646835f
C1257 a_n22294_n2937# dvss 0.502711f
C1258 a_n22672_n10337# dvss 0.639742f
C1259 a_n23050_n2937# dvss 0.502711f
C1260 a_n23428_n10337# dvss 0.639742f
C1261 a_n23806_n2937# dvss 0.502711f
C1262 a_n24184_n10337# dvss 0.639742f
C1263 a_n24562_n2937# dvss 0.502711f
C1264 a_n24940_n10337# dvss 0.639742f
C1265 a_n25318_n2937# dvss 0.502711f
C1266 a_n25696_n10337# dvss 0.639742f
C1267 a_n26074_n2937# dvss 0.502711f
C1268 a_n26452_n10337# dvss 0.639742f
C1269 a_n26830_n2937# dvss 0.502711f
C1270 a_n27208_n10337# dvss 0.614478f
C1271 ibias_gen_0.isrc_sel_b dvss 1.33811f
C1272 ibias_gen_0.isrc_sel dvss 5.28446f
C1273 ibias_gen_0.ena_b dvss 1.24326f
C1274 comparator_0.ibias dvss 2.77043f
C1275 ibias_gen_0.vp1 dvss 4.798203f
C1276 schmitt_trigger_0.in dvss 0.409716p
C1277 a_n8195_9395# dvss 0.502711f
C1278 a_n8573_1995# dvss 0.502711f
C1279 a_n8951_9395# dvss 0.502711f
C1280 a_n9329_1995# dvss 0.502711f
C1281 a_n9707_9395# dvss 0.502711f
C1282 a_n10085_1995# dvss 0.502711f
C1283 a_n10463_9395# dvss 0.502711f
C1284 a_n10841_1995# dvss 0.502711f
C1285 a_n11219_9395# dvss 0.502711f
C1286 a_n11597_1995# dvss 0.502711f
C1287 a_n11975_9395# dvss 0.502711f
C1288 a_n12353_1995# dvss 0.502711f
C1289 a_n12731_9395# dvss 0.502711f
C1290 a_n13109_1995# dvss 0.502711f
C1291 a_n13487_9395# dvss 0.502711f
C1292 a_n13865_1995# dvss 0.502711f
C1293 a_n14243_9395# dvss 0.502711f
C1294 a_n14621_1995# dvss 0.502711f
C1295 vl dvss 7.14205f
C1296 a_n14999_9395# dvss 0.502711f
C1297 dcomp3v3 dvss 1.22649f
C1298 comparator_1.n1 dvss 1.35962f
C1299 comparator_1.n0 dvss 0.750897f
C1300 comparator_1.vm dvss 4.47408f
C1301 comparator_1.vn dvss 4.961259f
C1302 ibias_gen_0.ibias0 dvss 0.517421f
C1303 comparator_1.ena_b dvss 0.625987f
C1304 comparator_0.ena dvss 9.82006f
C1305 comparator_1.vnn dvss 30.1825f
C1306 comparator_1.vpp dvss 29.323698f
C1307 comparator_0.vt dvss 11.7607f
C1308 comparator_1.vt dvss 4.36096f
C1309 rstring_mux_0.vtrip0.t0 dvss 0.791904f
C1310 rstring_mux_0.vtrip0.n0 dvss 0.190942f
C1311 rstring_mux_0.vtrip0.n1 dvss 0.125183f
C1312 rstring_mux_0.vtrip0.n2 dvss 0.776085f
C1313 rstring_mux_0.vtrip0.n3 dvss 0.190927f
C1314 rstring_mux_0.vtrip0.n4 dvss 0.125183f
C1315 rstring_mux_0.vtrip0.n5 dvss 1.22742f
C1316 rstring_mux_0.vtrip0.n6 dvss 2.02058f
C1317 rstring_mux_0.vtrip0.n7 dvss 1.79541f
C1318 rstring_mux_0.vtrip0.t5 dvss 0.169825f
C1319 ibias_gen_0.ve.n0 dvss -11.7115f
C1320 ibias_gen_0.ve.t1 dvss 11.8608f
C1321 ibias_gen_0.ve.t2 dvss 0.116976f
C1322 ibias_gen_0.ve.t3 dvss 0.116976f
C1323 ibias_gen_0.ve.n2 dvss 0.462255f
C1324 ibias_gen_0.ve.t4 dvss 0.116976f
C1325 ibias_gen_0.ve.t0 dvss 0.116976f
C1326 ibias_gen_0.ve.n3 dvss 0.496159f
C1327 ibias_gen_0.ve.n4 dvss 9.54037f
C1328 ibias_gen_0.ve.n5 dvss 10.730499f
C1329 rstring_mux_0.vtrip6.t5 dvss 0.172669f
C1330 rstring_mux_0.vtrip6.n0 dvss 0.187027f
C1331 rstring_mux_0.vtrip6.n1 dvss 0.122626f
C1332 rstring_mux_0.vtrip6.n2 dvss 0.800766f
C1333 rstring_mux_0.vtrip6.n3 dvss 0.187027f
C1334 rstring_mux_0.vtrip6.n4 dvss 0.122626f
C1335 rstring_mux_0.vtrip6.n5 dvss 1.249f
C1336 rstring_mux_0.vtrip6.n6 dvss 1.9489f
C1337 rstring_mux_0.vtrip6.n7 dvss 2.19091f
C1338 rstring_mux_0.vtrip6.t0 dvss 0.733177f
C1339 rstring_mux_0.vtrip1.t7 dvss 0.216167f
C1340 rstring_mux_0.vtrip1.n0 dvss 0.234604f
C1341 rstring_mux_0.vtrip1.n1 dvss 0.15382f
C1342 rstring_mux_0.vtrip1.n2 dvss 0.961398f
C1343 rstring_mux_0.vtrip1.n3 dvss 0.234604f
C1344 rstring_mux_0.vtrip1.n4 dvss 0.15382f
C1345 rstring_mux_0.vtrip1.n5 dvss 1.52407f
C1346 rstring_mux_0.vtrip1.n6 dvss 1.30427f
C1347 rstring_mux_0.vtrip1.n7 dvss 3.51872f
C1348 rstring_mux_0.vtrip1.t0 dvss 0.21619f
C1349 rstring_mux_0.vtrip5.t9 dvss 0.169149f
C1350 rstring_mux_0.vtrip5.n0 dvss 0.183575f
C1351 rstring_mux_0.vtrip5.n1 dvss 0.120363f
C1352 rstring_mux_0.vtrip5.n2 dvss 1.20735f
C1353 rstring_mux_0.vtrip5.n3 dvss 0.183575f
C1354 rstring_mux_0.vtrip5.n4 dvss 0.120363f
C1355 rstring_mux_0.vtrip5.n5 dvss 0.742428f
C1356 rstring_mux_0.vtrip5.n6 dvss 0.936052f
C1357 rstring_mux_0.vtrip5.n7 dvss 2.7123f
C1358 rstring_mux_0.vtrip5.t8 dvss 0.169167f
C1359 schmitt_trigger_0.out.n5 dvss 0.689226f
C1360 schmitt_trigger_0.out.t11 dvss 0.155689f
C1361 schmitt_trigger_0.out.t5 dvss 0.155538f
C1362 schmitt_trigger_0.out.n6 dvss 0.163942f
C1363 schmitt_trigger_0.out.t4 dvss 0.155622f
C1364 schmitt_trigger_0.out.n7 dvss 0.113412f
C1365 schmitt_trigger_0.out.t12 dvss 0.162392f
C1366 schmitt_trigger_0.out.n8 dvss 0.688643f
C1367 schmitt_trigger_0.out.n9 dvss 0.41845f
C1368 schmitt_trigger_0.out.n10 dvss 0.606738f
C1369 schmitt_trigger_0.out.n11 dvss 0.342028f
C1370 ibias_gen_0.vstart.n0 dvss 1.41043f
C1371 ibias_gen_0.vstart.n1 dvss 0.258324f
C1372 ibias_gen_0.vstart.t0 dvss 0.344828f
C1373 ibias_gen_0.vstart.n2 dvss 0.255572f
C1374 ibias_gen_0.vstart.n3 dvss 0.260069f
C1375 ibias_gen_0.vstart.n4 dvss 0.255572f
C1376 ibias_gen_0.vstart.n5 dvss 0.750761f
C1377 ibias_gen_0.vstart.n6 dvss 0.398642f
C1378 ibias_gen_0.vstart.n7 dvss 0.255572f
C1379 rstring_mux_0.vtrip3.t9 dvss 0.157727f
C1380 rstring_mux_0.vtrip3.n0 dvss 0.17118f
C1381 rstring_mux_0.vtrip3.n1 dvss 0.112235f
C1382 rstring_mux_0.vtrip3.n2 dvss 0.753957f
C1383 rstring_mux_0.vtrip3.n3 dvss 0.17118f
C1384 rstring_mux_0.vtrip3.n4 dvss 0.112235f
C1385 rstring_mux_0.vtrip3.n5 dvss 1.08769f
C1386 rstring_mux_0.vtrip3.n6 dvss 0.877189f
C1387 rstring_mux_0.vtrip3.n7 dvss 2.47396f
C1388 rstring_mux_0.vtrip3.t0 dvss 0.157744f
C1389 ibias_gen_0.vn1.n0 dvss 0.745323f
C1390 ibias_gen_0.vn1.t1 dvss 2.11164f
C1391 ibias_gen_0.vn1.t15 dvss 2.11164f
C1392 ibias_gen_0.vn1.t10 dvss 2.19722f
C1393 ibias_gen_0.vn1.n2 dvss 1.40052f
C1394 ibias_gen_0.vn1.t17 dvss 2.11164f
C1395 ibias_gen_0.vn1.t14 dvss 2.19722f
C1396 ibias_gen_0.vn1.n3 dvss 1.3685f
C1397 ibias_gen_0.vn1.n4 dvss 0.140807f
C1398 ibias_gen_0.vn1.t11 dvss 2.11164f
C1399 ibias_gen_0.vn1.t12 dvss 2.19722f
C1400 ibias_gen_0.vn1.n5 dvss 1.40052f
C1401 ibias_gen_0.vn1.t13 dvss 2.11164f
C1402 ibias_gen_0.vn1.t16 dvss 2.19722f
C1403 ibias_gen_0.vn1.n6 dvss 1.3685f
C1404 ibias_gen_0.vn1.n7 dvss 0.140807f
C1405 ibias_gen_0.vn1.n8 dvss 0.110984f
C1406 ibias_gen_0.vn1.n9 dvss 0.705651f
C1407 ibias_gen_0.vn1.t3 dvss 2.15704f
C1408 ibias_gen_0.vn1.n10 dvss 0.71883f
C1409 ibias_gen_0.vn1.n12 dvss 0.218051f
C1410 ibias_gen_0.vn1.n13 dvss 0.120433f
C1411 ibias_gen_0.vp1.n0 dvss 2.2551f
C1412 ibias_gen_0.vp1.t6 dvss 2.72493f
C1413 ibias_gen_0.vp1.n1 dvss 0.130918f
C1414 ibias_gen_0.vp1.n2 dvss 0.257085f
C1415 ibias_gen_0.vp1.n3 dvss 2.14115f
C1416 ibias_gen_0.vp1.t8 dvss 2.72114f
C1417 ibias_gen_0.vp1.n4 dvss 0.225585f
C1418 ibias_gen_0.vp1.n5 dvss 0.978301f
C1419 ibias_gen_0.vp1.n6 dvss 0.154917f
C1420 ibias_gen_0.vp1.n7 dvss 0.213443f
C1421 ibias_gen_0.vp1.n8 dvss 0.168888f
C1422 ibias_gen_0.vp1.n9 dvss 0.998605f
C1423 ibias_gen_0.vp1.n10 dvss 0.168888f
C1424 ibias_gen_0.vp1.n11 dvss 0.677866f
C1425 ibias_gen_0.vp1.n12 dvss 0.163248f
C1426 ibias_gen_0.vp1.n13 dvss 0.666034f
C1427 ibias_gen_0.vp1.n14 dvss 0.19773f
C1428 ibias_gen_0.vp1.n15 dvss 0.829697f
C1429 rstring_mux_0.vtrip2.t3 dvss 0.211519f
C1430 rstring_mux_0.vtrip2.n0 dvss 0.229108f
C1431 rstring_mux_0.vtrip2.n1 dvss 0.150216f
C1432 rstring_mux_0.vtrip2.n2 dvss 0.947831f
C1433 rstring_mux_0.vtrip2.n3 dvss 0.229108f
C1434 rstring_mux_0.vtrip2.n4 dvss 0.150216f
C1435 rstring_mux_0.vtrip2.n5 dvss 1.50485f
C1436 rstring_mux_0.vtrip2.n6 dvss 2.43692f
C1437 rstring_mux_0.vtrip2.n7 dvss 2.81264f
C1438 rstring_mux_0.vtrip2.t2 dvss 0.898141f
C1439 rstring_mux_0.vtrip7.t1 dvss 0.16069f
C1440 rstring_mux_0.vtrip7.n0 dvss 0.174395f
C1441 rstring_mux_0.vtrip7.n1 dvss 0.114343f
C1442 rstring_mux_0.vtrip7.n2 dvss 0.752155f
C1443 rstring_mux_0.vtrip7.n3 dvss 0.174395f
C1444 rstring_mux_0.vtrip7.n4 dvss 0.114343f
C1445 rstring_mux_0.vtrip7.n5 dvss 1.19247f
C1446 rstring_mux_0.vtrip7.n6 dvss 0.918289f
C1447 rstring_mux_0.vtrip7.n7 dvss 2.50533f
C1448 rstring_mux_0.vtrip7.t0 dvss 0.160707f
C1449 ibias_gen_0.vp.n0 dvss 0.431943f
C1450 ibias_gen_0.vp.t4 dvss 0.188332f
C1451 ibias_gen_0.vp.n3 dvss 0.662608f
C1452 ibias_gen_0.vp.t11 dvss 1.71268f
C1453 ibias_gen_0.vp.n4 dvss 1.29098f
C1454 ibias_gen_0.vp.t8 dvss 1.65245f
C1455 ibias_gen_0.vp.n5 dvss 1.29098f
C1456 ibias_gen_0.vp.t7 dvss 1.65245f
C1457 ibias_gen_0.vp.n6 dvss 1.29098f
C1458 ibias_gen_0.vp.t9 dvss 1.68256f
C1459 ibias_gen_0.vp.n7 dvss 0.597984f
C1460 ibias_gen_0.vp.t10 dvss 2.31092f
C1461 ibias_gen_0.vp.t12 dvss 2.34104f
C1462 ibias_gen_0.vp.n8 dvss 0.730243f
C1463 ibias_gen_0.vp.n9 dvss 1.1851f
C1464 ibias_gen_0.vp.n10 dvss 0.917156f
C1465 ibias_gen_0.vp.n12 dvss 0.488746f
C1466 ibias_gen_0.vr.n0 dvss 0.183081f
C1467 ibias_gen_0.vr.n1 dvss 0.161866f
C1468 ibias_gen_0.vr.n2 dvss 1.54735f
C1469 ibias_gen_0.vr.t4 dvss 0.540543f
C1470 ibias_gen_0.vp0.n0 dvss 0.777153f
C1471 ibias_gen_0.vp0.n1 dvss 0.217103f
C1472 ibias_gen_0.vp0.n3 dvss 0.886385f
C1473 ibias_gen_0.vp0.n5 dvss 0.157271f
C1474 ibias_gen_0.vp0.t8 dvss 1.72871f
C1475 ibias_gen_0.vp0.n6 dvss 1.47471f
C1476 ibias_gen_0.vp0.n7 dvss 0.724776f
C1477 ibias_gen_0.vp0.t13 dvss 1.76142f
C1478 ibias_gen_0.vp0.t12 dvss 1.69947f
C1479 ibias_gen_0.vp0.n8 dvss 1.47471f
C1480 ibias_gen_0.vp0.n9 dvss 0.800719f
C1481 ibias_gen_0.vp0.t10 dvss 1.69947f
C1482 ibias_gen_0.vp0.n10 dvss 0.798648f
C1483 ibias_gen_0.vp0.n11 dvss 0.128094f
C1484 ibias_gen_0.vp0.n12 dvss 0.98287f
C1485 ibias_gen_0.vp0.n13 dvss 1.07524f
C1486 ibias_gen_0.vp0.n14 dvss 0.139118f
C1487 ibias_gen_0.Mt4 dvss 1.25878f
C1488 ibias_gen_0.vn0.n0 dvss 0.935654f
C1489 ibias_gen_0.vn0.n1 dvss 1.39652f
C1490 ibias_gen_0.vn0.n2 dvss 0.142325f
C1491 ibias_gen_0.vn0.n3 dvss 0.874872f
C1492 ibias_gen_0.vn0.t19 dvss 2.24075f
C1493 ibias_gen_0.vn0.t3 dvss 2.19836f
C1494 ibias_gen_0.vn0.n4 dvss 0.920525f
C1495 ibias_gen_0.vn0.n5 dvss 0.111014f
C1496 ibias_gen_0.vn0.n6 dvss 0.198283f
C1497 ibias_gen_0.vn0.n7 dvss 0.161371f
C1498 ibias_gen_0.vn0.t1 dvss 2.16084f
C1499 ibias_gen_0.vn0.n8 dvss 1.01955f
C1500 ibias_gen_0.vn0.n9 dvss 1.87632f
C1501 ibias_gen_0.vn0.t20 dvss 2.16084f
C1502 ibias_gen_0.vn0.n10 dvss 1.71213f
C1503 ibias_gen_0.vn0.n11 dvss 0.975041f
C1504 ibias_gen_0.vn0.t9 dvss 0.202556f
C1505 ibias_gen_0.vn0.n12 dvss 0.12274f
C1506 ibias_gen_0.vn0.n13 dvss 0.12274f
C1507 ibias_gen_0.vn0.n14 dvss 0.12274f
C1508 ibias_gen_0.vn0.n15 dvss 0.12274f
C1509 ibias_gen_0.vn0.n16 dvss 0.12274f
C1510 vbg_1v2.n0 dvss 0.938703f
C1511 vbg_1v2.t21 dvss 1.50218f
C1512 vbg_1v2.t33 dvss 1.37455f
C1513 vbg_1v2.n1 dvss 0.934892f
C1514 vbg_1v2.t28 dvss 1.50218f
C1515 vbg_1v2.n4 dvss 0.934892f
C1516 vbg_1v2.t0 dvss 1.37455f
C1517 vbg_1v2.n5 dvss 0.934892f
C1518 vbg_1v2.t2 dvss 1.50218f
C1519 vbg_1v2.n8 dvss 0.934892f
C1520 vbg_1v2.t10 dvss 1.37455f
C1521 vbg_1v2.n9 dvss 0.934892f
C1522 vbg_1v2.t18 dvss 1.50218f
C1523 vbg_1v2.n12 dvss 0.934892f
C1524 vbg_1v2.t31 dvss 1.37455f
C1525 vbg_1v2.n13 dvss 0.934892f
C1526 vbg_1v2.t1 dvss 1.50218f
C1527 vbg_1v2.n16 dvss 0.934892f
C1528 vbg_1v2.t9 dvss 1.37455f
C1529 vbg_1v2.n17 dvss 0.934892f
C1530 vbg_1v2.t17 dvss 1.50218f
C1531 vbg_1v2.n20 dvss 0.934892f
C1532 vbg_1v2.t29 dvss 1.37455f
C1533 vbg_1v2.n21 dvss 0.934892f
C1534 vbg_1v2.t25 dvss 1.50218f
C1535 vbg_1v2.n24 dvss 0.934892f
C1536 vbg_1v2.t37 dvss 1.37455f
C1537 vbg_1v2.n25 dvss 0.934892f
C1538 vbg_1v2.t40 dvss 1.50218f
C1539 vbg_1v2.n28 dvss 0.934892f
C1540 vbg_1v2.t6 dvss 1.37455f
C1541 vbg_1v2.n29 dvss 0.934892f
C1542 vbg_1v2.n30 dvss 0.740506f
C1543 vbg_1v2.n31 dvss 0.938703f
C1544 vbg_1v2.t19 dvss 1.50218f
C1545 vbg_1v2.t35 dvss 1.37455f
C1546 vbg_1v2.n32 dvss 0.934892f
C1547 vbg_1v2.t11 dvss 1.50218f
C1548 vbg_1v2.n35 dvss 0.934892f
C1549 vbg_1v2.t26 dvss 1.37455f
C1550 vbg_1v2.n36 dvss 0.934892f
C1551 vbg_1v2.t36 dvss 1.50218f
C1552 vbg_1v2.n39 dvss 0.934892f
C1553 vbg_1v2.t7 dvss 1.37455f
C1554 vbg_1v2.n40 dvss 0.934892f
C1555 vbg_1v2.t23 dvss 1.50218f
C1556 vbg_1v2.n43 dvss 0.934892f
C1557 vbg_1v2.t38 dvss 1.37455f
C1558 vbg_1v2.n44 dvss 0.934892f
C1559 vbg_1v2.t4 dvss 1.50218f
C1560 vbg_1v2.n47 dvss 0.934892f
C1561 vbg_1v2.t16 dvss 1.37455f
C1562 vbg_1v2.n48 dvss 0.934892f
C1563 vbg_1v2.t24 dvss 1.50218f
C1564 vbg_1v2.n51 dvss 0.934892f
C1565 vbg_1v2.t39 dvss 1.37455f
C1566 vbg_1v2.n52 dvss 0.934892f
C1567 vbg_1v2.t14 dvss 1.50218f
C1568 vbg_1v2.n55 dvss 0.934892f
C1569 vbg_1v2.t32 dvss 1.37455f
C1570 vbg_1v2.n56 dvss 0.934892f
C1571 vbg_1v2.t12 dvss 1.50218f
C1572 vbg_1v2.n59 dvss 0.934892f
C1573 vbg_1v2.t27 dvss 1.37455f
C1574 vbg_1v2.n60 dvss 0.934892f
C1575 vbg_1v2.n61 dvss 1.17468f
C1576 vbg_1v2.n62 dvss 1.48365f
C1577 vbg_1v2.t34 dvss 0.2708f
C1578 vbg_1v2.n67 dvss 0.182117f
C1579 vbg_1v2.t30 dvss 0.270576f
C1580 vbg_1v2.n68 dvss 0.182117f
C1581 vbg_1v2.t20 dvss 0.270576f
C1582 vbg_1v2.t15 dvss 0.270576f
C1583 vbg_1v2.t8 dvss 0.270576f
C1584 vbg_1v2.t5 dvss 0.270576f
C1585 vbg_1v2.t3 dvss 0.270576f
C1586 vbg_1v2.t41 dvss 0.270576f
C1587 vbg_1v2.t13 dvss 0.270576f
C1588 vbg_1v2.t22 dvss 0.270576f
C1589 schmitt_trigger_0.m.n2 dvss 0.65613f
C1590 schmitt_trigger_0.m.n4 dvss 0.195435f
C1591 schmitt_trigger_0.m.t17 dvss 0.161114f
C1592 schmitt_trigger_0.m.t15 dvss 0.164304f
C1593 schmitt_trigger_0.m.t14 dvss 0.16415f
C1594 schmitt_trigger_0.m.n5 dvss 0.16975f
C1595 schmitt_trigger_0.m.t16 dvss 0.16428f
C1596 schmitt_trigger_0.m.n6 dvss 0.3748f
C1597 schmitt_trigger_0.m.n7 dvss 0.537335f
C1598 schmitt_trigger_0.m.n10 dvss 0.732652f
C1599 schmitt_trigger_0.m.n11 dvss 0.312554f
C1600 schmitt_trigger_0.m.n13 dvss 0.192206f
C1601 schmitt_trigger_0.m.n15 dvss 0.222965f
C1602 schmitt_trigger_0.in.t7 dvss 2.34931f
C1603 schmitt_trigger_0.in.t14 dvss 1.26511f
C1604 schmitt_trigger_0.in.n5 dvss 1.42394f
C1605 schmitt_trigger_0.in.t12 dvss 1.26511f
C1606 schmitt_trigger_0.in.n6 dvss 1.2565f
C1607 schmitt_trigger_0.in.t6 dvss 1.26511f
C1608 schmitt_trigger_0.in.n7 dvss 1.2565f
C1609 schmitt_trigger_0.in.t13 dvss 1.26511f
C1610 schmitt_trigger_0.in.n8 dvss 1.2565f
C1611 schmitt_trigger_0.in.t11 dvss 1.26511f
C1612 schmitt_trigger_0.in.n9 dvss 1.34081f
C1613 rstring_mux_0.vtop.n0 dvss 0.188061f
C1614 rstring_mux_0.vtop.n1 dvss 0.186982f
C1615 rstring_mux_0.vtop.n2 dvss 1.02937f
C1616 rstring_mux_0.vtop.n3 dvss 0.163921f
C1617 rstring_mux_0.vtop.n4 dvss 0.697228f
C1618 rstring_mux_0.vtop.n5 dvss 0.262825f
C1619 rstring_mux_0.vtop.n6 dvss 0.186982f
C1620 rstring_mux_0.vtop.n7 dvss 0.567273f
C1621 rstring_mux_0.vtop.n8 dvss 0.186982f
C1622 rstring_mux_0.vtop.n9 dvss 0.567273f
C1623 rstring_mux_0.vtop.n10 dvss 0.186982f
C1624 rstring_mux_0.vtop.n11 dvss 0.567273f
C1625 rstring_mux_0.vtop.n12 dvss 0.188542f
C1626 rstring_mux_0.vtop.n13 dvss 0.741617f
C1627 rstring_mux_0.vtop.n14 dvss 0.163921f
C1628 rstring_mux_0.vtop.n15 dvss 0.694975f
C1629 rstring_mux_0.vtop.t17 dvss 2.67225f
C1630 rc_osc_0.n.t11 dvss 0.143388f
C1631 rc_osc_0.n.t9 dvss 0.143249f
C1632 rc_osc_0.n.n2 dvss 0.164777f
C1633 rc_osc_0.n.t13 dvss 0.143249f
C1634 rc_osc_0.n.n3 dvss 0.156263f
C1635 rc_osc_0.n.t6 dvss 0.14446f
C1636 rc_osc_0.n.n4 dvss 0.529644f
C1637 rc_osc_0.n.t7 dvss 0.287357f
C1638 rc_osc_0.n.t12 dvss 0.286497f
C1639 rc_osc_0.n.n5 dvss 0.277287f
C1640 rc_osc_0.n.t8 dvss 0.287213f
C1641 rc_osc_0.n.n6 dvss 0.196012f
C1642 rc_osc_0.n.t10 dvss 0.283047f
C1643 rc_osc_0.n.n7 dvss 0.360416f
C1644 rc_osc_0.n.n8 dvss 0.222174f
C1645 rc_osc_0.n.n9 dvss 0.477653f
C1646 rc_osc_0.n.n10 dvss 0.555032f
C1647 dvdd.n184 dvss 0.149811f
C1648 dvdd.n204 dvss 0.108058f
C1649 dvdd.n205 dvss 0.108058f
C1650 dvdd.n209 dvss 0.107566f
C1651 dvdd.n210 dvss 0.126887f
C1652 dvdd.n267 dvss 0.691637f
C1653 dvdd.n268 dvss 0.202814f
C1654 dvdd.n269 dvss 0.440047f
C1655 dvdd.n270 dvss 0.439981f
C1656 dvdd.n271 dvss 1.65526f
C1657 dvdd.n272 dvss 0.441923f
C1658 dvdd.n273 dvss 1.68313f
C1659 dvdd.n274 dvss 1.655f
C1660 dvdd.n275 dvss 1.68287f
C1661 dvdd.n276 dvss 0.441856f
C1662 dvdd.n277 dvss 0.202783f
C1663 dvdd.n278 dvss 1.00601f
C1664 dvdd.n280 dvss 0.41383f
C1665 dvdd.n281 dvss 0.114124f
C1666 dvdd.n351 dvss 0.509148f
C1667 dvdd.n460 dvss 0.550925f
C1668 dvdd.n463 dvss 0.133555f
C1669 dvdd.n464 dvss 1.80993f
C1670 dvdd.n465 dvss 0.477551f
C1671 dvdd.n466 dvss 1.03683f
C1672 dvdd.n467 dvss 1.03683f
C1673 dvdd.n468 dvss 3.95208f
C1674 dvdd.n469 dvss 1.04032f
C1675 dvdd.n470 dvss 4.00553f
C1676 dvdd.n471 dvss 3.95208f
C1677 dvdd.n472 dvss 4.00553f
C1678 dvdd.n473 dvss 1.04032f
C1679 dvdd.n474 dvss 0.477551f
C1680 dvdd.n475 dvss 2.25176f
C1681 dvdd.n476 dvss 0.176366f
C1682 dvdd.n496 dvss 0.128459f
C1683 dvdd.n502 dvss 0.233225f
C1684 dvdd.t64 dvss 0.206708f
C1685 dvdd.t62 dvss 0.154382f
C1686 dvdd.t222 dvss 0.154382f
C1687 dvdd.t282 dvss 0.154382f
C1688 dvdd.t284 dvss 0.154382f
C1689 dvdd.t286 dvss 0.154382f
C1690 dvdd.t123 dvss 0.17881f
C1691 dvdd.t58 dvss 0.227665f
C1692 dvdd.t220 dvss 0.252092f
C1693 dvdd.t60 dvss 0.129466f
C1694 dvdd.n503 dvss 0.101618f
C1695 dvdd.t189 dvss 0.175389f
C1696 dvdd.t191 dvss 0.154382f
C1697 dvdd.t187 dvss 0.154382f
C1698 dvdd.t193 dvss 0.154382f
C1699 dvdd.t183 dvss 0.154382f
C1700 dvdd.t185 dvss 0.139237f
C1701 dvdd.t125 dvss 0.108946f
C1702 dvdd.t95 dvss 0.108946f
C1703 dvdd.t118 dvss 0.144122f
C1704 dvdd.t131 dvss 0.14852f
C1705 dvdd.t115 dvss 0.110901f
C1706 dvdd.t133 dvss 0.146909f
C1707 dvdd.n504 dvss 0.204598f
C1708 dvdd.n509 dvss 0.945498f
C1709 dvdd.n513 dvss 0.72682f
C1710 dvdd.n514 dvss 1.91741f
C1711 dvdd.n515 dvss 0.162528f
C1712 avdd.t153 dvss 1.97912f
C1713 avdd.t159 dvss 0.809969f
C1714 avdd.t14 dvss 1.32299f
C1715 avdd.t517 dvss 1.97912f
C1716 avdd.t519 dvss 0.809969f
C1717 avdd.t456 dvss 1.32299f
C1718 avdd.t454 dvss 1.97912f
C1719 avdd.t452 dvss 0.809969f
C1720 avdd.t209 dvss 1.32299f
C1721 avdd.t172 dvss 1.97912f
C1722 avdd.t584 dvss 0.809969f
C1723 avdd.t444 dvss 1.32299f
C1724 avdd.t406 dvss 1.97912f
C1725 avdd.t404 dvss 0.809969f
C1726 avdd.t484 dvss 1.32299f
C1727 avdd.t0 dvss 1.97912f
C1728 avdd.t120 dvss 0.809969f
C1729 avdd.t205 dvss 1.32299f
C1730 avdd.t515 dvss 1.97912f
C1731 avdd.t513 dvss 0.809969f
C1732 avdd.t414 dvss 1.32299f
C1733 avdd.t450 dvss 1.97912f
C1734 avdd.t486 dvss 0.809969f
C1735 avdd.t501 dvss 1.32299f
C1736 avdd.t52 dvss 0.265371f
C1737 avdd.n69 dvss 0.644224f
C1738 avdd.n73 dvss 0.14577f
C1739 avdd.n74 dvss 0.688565f
C1740 avdd.t165 dvss 1.39358f
C1741 avdd.n77 dvss 1.22533f
C1742 avdd.n87 dvss 0.223055f
C1743 avdd.n93 dvss 0.500334f
C1744 avdd.t565 dvss 0.265371f
C1745 avdd.n94 dvss 0.295778f
C1746 avdd.n95 dvss 0.425699f
C1747 avdd.n98 dvss 0.370413f
C1748 avdd.n99 dvss 0.530741f
C1749 avdd.t50 dvss 1.29921f
C1750 avdd.t421 dvss 0.237728f
C1751 avdd.n100 dvss 0.480984f
C1752 avdd.n118 dvss 0.223055f
C1753 avdd.n125 dvss 1.39126f
C1754 avdd.n128 dvss 1.18013f
C1755 avdd.n146 dvss 0.223055f
C1756 avdd.n153 dvss 1.39126f
C1757 avdd.n156 dvss 1.18013f
C1758 avdd.n174 dvss 0.223055f
C1759 avdd.n181 dvss 1.39126f
C1760 avdd.n184 dvss 1.18013f
C1761 avdd.n202 dvss 0.223055f
C1762 avdd.n209 dvss 1.39126f
C1763 avdd.n212 dvss 1.18013f
C1764 avdd.n230 dvss 0.223055f
C1765 avdd.n237 dvss 1.39126f
C1766 avdd.n240 dvss 1.18013f
C1767 avdd.n258 dvss 0.223055f
C1768 avdd.n265 dvss 1.39126f
C1769 avdd.n268 dvss 1.18013f
C1770 avdd.n286 dvss 0.223055f
C1771 avdd.n293 dvss 1.39126f
C1772 avdd.n296 dvss 1.18013f
C1773 avdd.n314 dvss 0.223055f
C1774 avdd.n321 dvss 1.39126f
C1775 avdd.n324 dvss 1.18013f
C1776 avdd.t215 dvss 1.97912f
C1777 avdd.t416 dvss 0.809969f
C1778 avdd.t16 dvss 1.32299f
C1779 avdd.t110 dvss 1.97912f
C1780 avdd.t496 dvss 0.809969f
C1781 avdd.t482 dvss 1.32299f
C1782 avdd.t442 dvss 1.97912f
C1783 avdd.t440 dvss 0.809969f
C1784 avdd.t410 dvss 1.32299f
C1785 avdd.t116 dvss 1.97912f
C1786 avdd.t535 dvss 0.809969f
C1787 avdd.t493 dvss 1.32299f
C1788 avdd.t112 dvss 1.97912f
C1789 avdd.t114 dvss 0.809969f
C1790 avdd.t4 dvss 1.32299f
C1791 avdd.t54 dvss 1.97912f
C1792 avdd.t56 dvss 0.809969f
C1793 avdd.t567 dvss 1.32299f
C1794 avdd.t528 dvss 1.97912f
C1795 avdd.t607 dvss 0.809969f
C1796 avdd.t224 dvss 1.32299f
C1797 avdd.t10 dvss 1.97912f
C1798 avdd.t12 dvss 0.809969f
C1799 avdd.t526 dvss 1.32299f
C1800 avdd.t8 dvss 0.265371f
C1801 avdd.n405 dvss 0.640917f
C1802 avdd.n409 dvss 0.14577f
C1803 avdd.n410 dvss 0.688565f
C1804 avdd.t48 dvss 1.39328f
C1805 avdd.n413 dvss 1.22533f
C1806 avdd.n423 dvss 0.223055f
C1807 avdd.n429 dvss 0.49757f
C1808 avdd.t221 dvss 0.265371f
C1809 avdd.n430 dvss 0.295778f
C1810 avdd.n431 dvss 0.425699f
C1811 avdd.n434 dvss 0.370413f
C1812 avdd.n435 dvss 0.530741f
C1813 avdd.t6 dvss 1.29921f
C1814 avdd.t102 dvss 0.237728f
C1815 avdd.n436 dvss 0.480984f
C1816 avdd.n454 dvss 0.223055f
C1817 avdd.n461 dvss 1.39126f
C1818 avdd.n464 dvss 1.18013f
C1819 avdd.n482 dvss 0.223055f
C1820 avdd.n489 dvss 1.39126f
C1821 avdd.n492 dvss 1.18013f
C1822 avdd.n510 dvss 0.223055f
C1823 avdd.n517 dvss 1.39126f
C1824 avdd.n520 dvss 1.18013f
C1825 avdd.n538 dvss 0.223055f
C1826 avdd.n545 dvss 1.39126f
C1827 avdd.n548 dvss 1.18013f
C1828 avdd.n566 dvss 0.223055f
C1829 avdd.n573 dvss 1.39126f
C1830 avdd.n576 dvss 1.18013f
C1831 avdd.n594 dvss 0.223055f
C1832 avdd.n601 dvss 1.39126f
C1833 avdd.n604 dvss 1.18013f
C1834 avdd.n622 dvss 0.223055f
C1835 avdd.n629 dvss 1.39126f
C1836 avdd.n632 dvss 1.18013f
C1837 avdd.n650 dvss 0.223055f
C1838 avdd.n657 dvss 1.39126f
C1839 avdd.n660 dvss 1.18013f
C1840 avdd.n672 dvss 4.69798f
C1841 avdd.n673 dvss 5.99918f
C1842 avdd.n674 dvss 5.24583f
C1843 avdd.t541 dvss 1.00017f
C1844 avdd.n680 dvss 0.592751f
C1845 avdd.n686 dvss 0.305482f
C1846 avdd.n687 dvss 0.115502f
C1847 avdd.n688 dvss 1.08469f
C1848 avdd.t253 dvss 0.777238f
C1849 avdd.n689 dvss 0.482557f
C1850 avdd.n690 dvss 1.06438f
C1851 avdd.n691 dvss 0.63618f
C1852 avdd.n692 dvss 2.09927f
C1853 avdd.n693 dvss 2.09927f
C1854 avdd.n694 dvss 0.63618f
C1855 avdd.n695 dvss 1.06488f
C1856 avdd.n697 dvss 0.315222f
C1857 avdd.t563 dvss 0.499357f
C1858 avdd.n704 dvss 0.187737f
C1859 avdd.n705 dvss 0.830596f
C1860 avdd.n706 dvss 0.824907f
C1861 avdd.t46 dvss 0.182048f
C1862 avdd.t408 dvss 0.182048f
C1863 avdd.n715 dvss 0.305482f
C1864 avdd.n717 dvss 0.210493f
C1865 avdd.n723 dvss 0.187737f
C1866 avdd.n725 dvss 0.830596f
C1867 avdd.n726 dvss 0.824907f
C1868 avdd.t157 dvss 0.182048f
C1869 avdd.t577 dvss 0.182048f
C1870 avdd.n735 dvss 0.305482f
C1871 avdd.n737 dvss 0.210493f
C1872 avdd.n743 dvss 0.187737f
C1873 avdd.n745 dvss 0.830596f
C1874 avdd.n746 dvss 0.824907f
C1875 avdd.t609 dvss 0.182048f
C1876 avdd.t207 dvss 0.182048f
C1877 avdd.n755 dvss 0.305482f
C1878 avdd.n757 dvss 0.210493f
C1879 avdd.n763 dvss 0.187737f
C1880 avdd.n765 dvss 0.830596f
C1881 avdd.n766 dvss 0.824907f
C1882 avdd.t579 dvss 0.182048f
C1883 avdd.t581 dvss 0.182048f
C1884 avdd.n775 dvss 0.305482f
C1885 avdd.n777 dvss 0.210493f
C1886 avdd.n783 dvss 0.187737f
C1887 avdd.n785 dvss 0.830596f
C1888 avdd.n786 dvss 0.824907f
C1889 avdd.t211 dvss 0.182048f
C1890 avdd.t532 dvss 0.651705f
C1891 avdd.n795 dvss 0.305482f
C1892 avdd.n797 dvss 0.210493f
C1893 avdd.n798 dvss 0.220841f
C1894 avdd.n799 dvss 0.159266f
C1895 avdd.n802 dvss 0.305482f
C1896 avdd.n808 dvss 0.824907f
C1897 avdd.n809 dvss 0.830596f
C1898 avdd.n810 dvss 0.187737f
C1899 avdd.n814 dvss 0.210493f
C1900 avdd.n815 dvss 0.305482f
C1901 avdd.n820 dvss 0.830596f
C1902 avdd.n821 dvss 0.187737f
C1903 avdd.t106 dvss 0.182048f
C1904 avdd.n822 dvss 0.824907f
C1905 avdd.n825 dvss 0.210493f
C1906 avdd.n827 dvss 0.305482f
C1907 avdd.n833 dvss 0.824907f
C1908 avdd.n834 dvss 0.830596f
C1909 avdd.n835 dvss 0.187737f
C1910 avdd.n839 dvss 0.210493f
C1911 avdd.n840 dvss 0.305482f
C1912 avdd.n845 dvss 0.830596f
C1913 avdd.n846 dvss 0.187737f
C1914 avdd.t118 dvss 0.182048f
C1915 avdd.n847 dvss 0.824907f
C1916 avdd.n850 dvss 0.210493f
C1917 avdd.n852 dvss 0.305482f
C1918 avdd.n858 dvss 0.824907f
C1919 avdd.n859 dvss 0.830596f
C1920 avdd.n860 dvss 0.187737f
C1921 avdd.n864 dvss 0.210493f
C1922 avdd.n865 dvss 0.305482f
C1923 avdd.n870 dvss 0.830596f
C1924 avdd.n871 dvss 0.187737f
C1925 avdd.t539 dvss 0.182048f
C1926 avdd.n872 dvss 0.824907f
C1927 avdd.n875 dvss 0.210493f
C1928 avdd.n877 dvss 0.305482f
C1929 avdd.n883 dvss 0.824907f
C1930 avdd.n884 dvss 0.830596f
C1931 avdd.n885 dvss 0.187737f
C1932 avdd.n889 dvss 0.210493f
C1933 avdd.n890 dvss 0.305482f
C1934 avdd.n895 dvss 0.830596f
C1935 avdd.n896 dvss 0.187737f
C1936 avdd.t104 dvss 0.182048f
C1937 avdd.n897 dvss 0.824907f
C1938 avdd.n900 dvss 0.210493f
C1939 avdd.n902 dvss 0.305482f
C1940 avdd.n908 dvss 0.824907f
C1941 avdd.n909 dvss 0.830596f
C1942 avdd.n910 dvss 0.187737f
C1943 avdd.n914 dvss 0.210493f
C1944 avdd.n915 dvss 0.305482f
C1945 avdd.n920 dvss 0.830596f
C1946 avdd.n921 dvss 0.187737f
C1947 avdd.t530 dvss 0.182048f
C1948 avdd.n922 dvss 0.824907f
C1949 avdd.n925 dvss 0.210493f
C1950 avdd.n926 dvss 0.305482f
C1951 avdd.n932 dvss 1.03262f
C1952 avdd.t309 dvss 0.777238f
C1953 avdd.t248 dvss 0.777238f
C1954 avdd.t338 dvss 0.777238f
C1955 avdd.t280 dvss 0.777238f
C1956 avdd.t380 dvss 0.777238f
C1957 avdd.t267 dvss 0.777238f
C1958 avdd.t398 dvss 0.777238f
C1959 avdd.t386 dvss 0.777238f
C1960 avdd.t373 dvss 0.777238f
C1961 avdd.t384 dvss 0.777238f
C1962 avdd.t302 dvss 0.777238f
C1963 avdd.t396 dvss 0.777238f
C1964 avdd.t400 dvss 0.777238f
C1965 avdd.t362 dvss 0.777238f
C1966 avdd.n933 dvss 0.483826f
C1967 avdd.n934 dvss 0.483826f
C1968 avdd.n935 dvss 0.483826f
C1969 avdd.n936 dvss 0.483826f
C1970 avdd.n937 dvss 0.483826f
C1971 avdd.n938 dvss 0.483826f
C1972 avdd.n939 dvss 0.377646f
C1973 avdd.n940 dvss 0.112949f
C1974 avdd.n941 dvss 0.477057f
C1975 avdd.n942 dvss 0.483826f
C1976 avdd.n943 dvss 0.483826f
C1977 avdd.n944 dvss 0.483826f
C1978 avdd.n945 dvss 0.483826f
C1979 avdd.n946 dvss 0.483826f
C1980 avdd.n947 dvss 0.496916f
C1981 avdd.n948 dvss 0.307641f
C1982 avdd.n949 dvss 2.49277f
C1983 avdd.n950 dvss 9.57984f
C1984 avdd.n951 dvss 0.822354f
C1985 avdd.n952 dvss 2.72536f
C1986 avdd.t226 dvss 2.86945f
C1987 avdd.n953 dvss 1.3892f
C1988 avdd.n954 dvss 0.213133f
C1989 avdd.n955 dvss 0.640478f
C1990 avdd.n956 dvss 0.190327f
C1991 avdd.n957 dvss 1.34232f
C1992 avdd.n958 dvss 1.42497f
C1993 avdd.n959 dvss 2.26261f
C1994 avdd.t227 dvss 48.5178f
C1995 avdd.n960 dvss 0.563898f
C1996 avdd.n961 dvss 2.71162f
C1997 avdd.n962 dvss 2.49618f
C1998 avdd.n963 dvss 1.54067f
C1999 avdd.n964 dvss 1.46547f
C2000 avdd.n965 dvss 0.197642f
C2001 avdd.n966 dvss 0.264953f
C2002 avdd.n967 dvss 0.449492f
C2003 avdd.n968 dvss 0.154989f
C2004 avdd.n969 dvss 0.16721f
C2005 avdd.t549 dvss 1.33689f
C2006 avdd.t174 dvss 1.85021f
C2007 avdd.n970 dvss 1.63778f
C2008 avdd.n971 dvss 0.449492f
C2009 avdd.t551 dvss 1.52228f
C2010 avdd.t543 dvss 1.67463f
C2011 avdd.n972 dvss 1.44258f
C2012 avdd.n973 dvss 0.16721f
C2013 avdd.n974 dvss 0.154989f
C2014 avdd.n975 dvss 0.123867f
C2015 avdd.n976 dvss 0.833717f
C2016 avdd.n977 dvss 2.1473f
C2017 avdd.n978 dvss 1.54067f
C2018 avdd.t22 dvss 46.0373f
C2019 avdd.t33 dvss 61.383f
C2020 avdd.t18 dvss 46.0373f
C2021 avdd.n979 dvss 1.42497f
C2022 avdd.n980 dvss 0.640478f
C2023 avdd.n982 dvss 0.258624f
C2024 avdd.n983 dvss 1.92926f
C2025 avdd.n984 dvss 1.78436f
C2026 avdd.n985 dvss 1.00681f
C2027 avdd.n987 dvss 0.460184f
C2028 avdd.n989 dvss 0.286865f
C2029 avdd.n991 dvss 0.286865f
C2030 avdd.n993 dvss 0.326308f
C2031 avdd.n995 dvss 0.326308f
C2032 avdd.n997 dvss 0.286865f
C2033 avdd.n999 dvss 0.286865f
C2034 avdd.n1001 dvss 0.286865f
C2035 avdd.n1003 dvss 0.286865f
C2036 avdd.n1005 dvss 0.286865f
C2037 avdd.n1007 dvss 0.258624f
C2038 avdd.n1008 dvss 0.115125f
C2039 avdd.n1010 dvss 0.247668f
C2040 avdd.n1011 dvss 2.57803f
C2041 avdd.n1012 dvss 0.880834f
C2042 avdd.n1013 dvss 0.978922f
C2043 avdd.n1014 dvss 0.993149f
C2044 avdd.n1015 dvss 4.22301f
C2045 avdd.n1016 dvss 4.22247f
C2046 avdd.n1017 dvss 15.931701f
C2047 avdd.n1018 dvss 1.02641f
C2048 avdd.n1019 dvss 0.99239f
C2049 avdd.n1020 dvss 0.901373f
C2050 avdd.n1021 dvss 1.80268f
C2051 avdd.n1022 dvss 0.880834f
C2052 avdd.n1023 dvss 1.53938f
C2053 avdd.n1024 dvss 0.115125f
C2054 avdd.n1025 dvss 0.142138f
C2055 avdd.n1026 dvss 0.136266f
C2056 avdd.n1027 dvss 0.127835f
C2057 avdd.n1028 dvss 0.78481f
C2058 avdd.n1029 dvss 2.8425f
C2059 avdd.n1030 dvss 3.13648f
C2060 avdd.n1031 dvss 2.83597f
C2061 avdd.n1032 dvss 0.794727f
C2062 avdd.n1033 dvss 0.166768f
C2063 avdd.n1034 dvss 0.236203f
C2064 avdd.t426 dvss 0.704956f
C2065 avdd.n1035 dvss 0.539054f
C2066 avdd.t436 dvss 0.704956f
C2067 avdd.t432 dvss 0.939941f
C2068 avdd.t434 dvss 0.939941f
C2069 avdd.t424 dvss 0.939941f
C2070 avdd.t430 dvss 1.1627f
C2071 avdd.n1036 dvss 1.5397f
C2072 avdd.t428 dvss 0.939941f
C2073 avdd.t438 dvss 0.939941f
C2074 avdd.t177 dvss 0.939941f
C2075 avdd.t175 dvss 1.1627f
C2076 avdd.n1037 dvss 1.5397f
C2077 avdd.n1038 dvss 0.18791f
C2078 avdd.n1039 dvss 0.172686f
C2079 avdd.n1040 dvss 0.317697f
C2080 avdd.n1041 dvss 0.172686f
C2081 avdd.n1043 dvss 0.286865f
C2082 avdd.n1045 dvss 0.286865f
C2083 avdd.n1047 dvss 0.286865f
C2084 avdd.n1049 dvss 0.286865f
C2085 avdd.n1051 dvss 0.286865f
C2086 avdd.n1053 dvss 0.326308f
C2087 avdd.n1055 dvss 0.326308f
C2088 avdd.n1057 dvss 0.286865f
C2089 avdd.n1059 dvss 0.286865f
C2090 avdd.n1061 dvss 0.460184f
C2091 avdd.n1062 dvss 3.62023f
C2092 avdd.n1063 dvss 2.72536f
C2093 avdd.n1064 dvss 0.170379f
C2094 avdd.n1065 dvss 0.326308f
C2095 avdd.t287 dvss 2.85263f
C2096 avdd.n1066 dvss 0.170379f
C2097 avdd.n1067 dvss 0.286865f
C2098 avdd.t382 dvss 2.85333f
C2099 avdd.n1068 dvss 0.170379f
C2100 avdd.t255 dvss 2.85333f
C2101 avdd.n1069 dvss 1.40632f
C2102 avdd.n1071 dvss 0.258624f
C2103 avdd.t391 dvss 2.85333f
C2104 avdd.n1072 dvss 1.40632f
C2105 avdd.n1074 dvss 0.286865f
C2106 avdd.n1075 dvss 0.286865f
C2107 avdd.t245 dvss 2.85333f
C2108 avdd.n1077 dvss 1.40632f
C2109 avdd.n1078 dvss 0.170379f
C2110 avdd.t375 dvss 2.85333f
C2111 avdd.n1080 dvss 1.40632f
C2112 avdd.n1081 dvss 0.170379f
C2113 avdd.n1082 dvss 0.170379f
C2114 avdd.n1083 dvss 1.40632f
C2115 avdd.n1085 dvss 0.286865f
C2116 avdd.t368 dvss 2.85333f
C2117 avdd.n1086 dvss 1.40632f
C2118 avdd.n1088 dvss 0.286865f
C2119 avdd.n1089 dvss 0.326308f
C2120 avdd.t366 dvss 2.85333f
C2121 avdd.n1091 dvss 1.40632f
C2122 avdd.n1092 dvss 0.209822f
C2123 avdd.t352 dvss 2.85263f
C2124 avdd.n1094 dvss 1.4013f
C2125 avdd.n1095 dvss 0.209822f
C2126 avdd.n1096 dvss 0.170379f
C2127 avdd.n1097 dvss 1.4013f
C2128 avdd.n1099 dvss 0.286865f
C2129 avdd.t289 dvss 2.85263f
C2130 avdd.n1100 dvss 1.4013f
C2131 avdd.n1102 dvss 0.286865f
C2132 avdd.n1103 dvss 0.460184f
C2133 avdd.t282 dvss 2.85263f
C2134 avdd.n1105 dvss 1.4013f
C2135 avdd.n1106 dvss 0.343698f
C2136 avdd.n1107 dvss 2.01084f
C2137 avdd.n1108 dvss 0.830753f
C2138 avdd.n1109 dvss 0.241516f
C2139 avdd.n1111 dvss 0.285283f
C2140 avdd.n1113 dvss 0.285283f
C2141 avdd.n1115 dvss 0.285283f
C2142 avdd.n1117 dvss 0.285283f
C2143 avdd.n1118 dvss 0.306627f
C2144 avdd.n1119 dvss 0.189145f
C2145 avdd.n1120 dvss 0.289183f
C2146 avdd.n1121 dvss 0.539054f
C2147 avdd.n1122 dvss 2.22853f
C2148 avdd.n1123 dvss 0.563898f
C2149 avdd.t25 dvss 61.383f
C2150 avdd.t246 dvss 48.5178f
C2151 avdd.n1124 dvss 0.834636f
C2152 avdd.n1125 dvss 1.42313f
C2153 avdd.n1126 dvss 19.5848f
C2154 avdd.n1127 dvss 1.19282f
C2155 avdd.n1128 dvss 0.713752f
C2156 avdd.n1129 dvss 0.217503f
C2157 avdd.n1130 dvss 0.247032f
C2158 avdd.n1131 dvss 0.115125f
C2159 avdd.n1132 dvss 0.213134f
C2160 avdd.t273 dvss 2.86945f
C2161 avdd.n1133 dvss 1.3892f
C2162 avdd.n1135 dvss 0.794824f
C2163 avdd.n1136 dvss 2.04908f
C2164 avdd.n1137 dvss 2.50608f
C2165 avdd.n1138 dvss 1.96847f
C2166 avdd.n1139 dvss 0.960954f
C2167 avdd.n1140 dvss 0.980125f
C2168 avdd.n1141 dvss 4.23964f
C2169 avdd.n1142 dvss 16.1996f
C2170 avdd.n1143 dvss 15.9296f
C2171 avdd.n1144 dvss 16.1996f
C2172 avdd.n1145 dvss 4.23964f
C2173 avdd.n1146 dvss 0.979544f
C2174 avdd.n1147 dvss 0.948763f
C2175 avdd.n1148 dvss 1.96847f
C2176 avdd.n1149 dvss 1.77298f
C2177 avdd.n1150 dvss 1.95878f
C2178 avdd.n1151 dvss 0.637456f
C2179 avdd.n1152 dvss 1.16091f
C2180 avdd.n1153 dvss 1.93485f
C2181 avdd.n1154 dvss 0.605048f
C2182 avdd.n1156 dvss 0.2402f
C2183 avdd.n1157 dvss 0.115125f
C2184 avdd.n1158 dvss 0.846056f
C2185 avdd.n1159 dvss 2.16083f
C2186 avdd.n1160 dvss 30.6915f
C2187 avdd.n1161 dvss 2.16083f
C2188 avdd.n1162 dvss 1.26669f
C2189 avdd.n1163 dvss 0.771102f
C2190 avdd.n1164 dvss 0.834636f
C2191 avdd.n1165 dvss 1.42313f
C2192 avdd.n1166 dvss 19.5848f
C2193 avdd.n1167 dvss 1.19282f
C2194 avdd.n1168 dvss 0.713752f
C2195 avdd.n1169 dvss 0.14348f
C2196 avdd.n1170 dvss 0.247032f
C2197 avdd.n1171 dvss 0.115125f
C2198 avdd.t393 dvss 2.85333f
C2199 avdd.n1172 dvss 1.40632f
C2200 avdd.n1173 dvss 0.142138f
C2201 avdd.t340 dvss 2.85333f
C2202 avdd.n1174 dvss 1.40632f
C2203 avdd.n1175 dvss 0.170379f
C2204 avdd.t388 dvss 2.85333f
C2205 avdd.n1176 dvss 1.40632f
C2206 avdd.n1177 dvss 0.170379f
C2207 avdd.t327 dvss 2.85333f
C2208 avdd.n1178 dvss 1.40632f
C2209 avdd.n1179 dvss 0.170379f
C2210 avdd.t332 dvss 2.85333f
C2211 avdd.n1180 dvss 1.40632f
C2212 avdd.n1181 dvss 0.170379f
C2213 avdd.t317 dvss 2.85333f
C2214 avdd.n1182 dvss 1.40632f
C2215 avdd.n1183 dvss 0.170379f
C2216 avdd.t314 dvss 2.85333f
C2217 avdd.n1184 dvss 1.40632f
C2218 avdd.n1185 dvss 0.209822f
C2219 avdd.t294 dvss 2.85263f
C2220 avdd.n1186 dvss 1.4013f
C2221 avdd.n1187 dvss 0.209822f
C2222 avdd.t257 dvss 2.85263f
C2223 avdd.n1188 dvss 1.4013f
C2224 avdd.n1189 dvss 0.170379f
C2225 avdd.t260 dvss 2.85263f
C2226 avdd.n1190 dvss 1.4013f
C2227 avdd.n1191 dvss 0.170379f
C2228 avdd.t250 dvss 2.85263f
C2229 avdd.n1192 dvss 1.4013f
C2230 avdd.n1193 dvss 0.343698f
C2231 avdd.n1194 dvss 1.32207f
C2232 avdd.n1195 dvss 0.516245f
C2233 avdd.n1196 dvss 1.04548f
C2234 avdd.n1197 dvss 0.774177f
C2235 avdd.n1198 dvss 2.72536f
C2236 avdd.t277 dvss 2.86945f
C2237 avdd.n1199 dvss 1.3892f
C2238 avdd.n1200 dvss 0.213133f
C2239 avdd.n1201 dvss 0.640478f
C2240 avdd.n1202 dvss 0.190327f
C2241 avdd.n1203 dvss 1.34232f
C2242 avdd.n1204 dvss 1.42497f
C2243 avdd.n1205 dvss 2.26261f
C2244 avdd.t236 dvss 48.5178f
C2245 avdd.n1206 dvss 0.563898f
C2246 avdd.n1207 dvss 2.71162f
C2247 avdd.n1208 dvss 2.49618f
C2248 avdd.n1209 dvss 1.54067f
C2249 avdd.n1210 dvss 1.46547f
C2250 avdd.n1211 dvss 0.197642f
C2251 avdd.n1212 dvss 0.264953f
C2252 avdd.n1213 dvss 0.449492f
C2253 avdd.n1214 dvss 0.154989f
C2254 avdd.n1215 dvss 0.16721f
C2255 avdd.t559 dvss 1.33689f
C2256 avdd.t524 dvss 1.85021f
C2257 avdd.n1216 dvss 1.63778f
C2258 avdd.n1217 dvss 0.449492f
C2259 avdd.t553 dvss 1.52228f
C2260 avdd.t561 dvss 1.67463f
C2261 avdd.n1218 dvss 1.44258f
C2262 avdd.n1219 dvss 0.16721f
C2263 avdd.n1220 dvss 0.154989f
C2264 avdd.n1221 dvss 0.123867f
C2265 avdd.n1222 dvss 0.833717f
C2266 avdd.n1223 dvss 2.1473f
C2267 avdd.n1224 dvss 1.54067f
C2268 avdd.t133 dvss 46.0373f
C2269 avdd.t123 dvss 61.383f
C2270 avdd.t125 dvss 46.0373f
C2271 avdd.n1225 dvss 1.42497f
C2272 avdd.n1226 dvss 0.640478f
C2273 avdd.n1228 dvss 0.258624f
C2274 avdd.n1229 dvss 1.92926f
C2275 avdd.n1230 dvss 1.78436f
C2276 avdd.n1231 dvss 1.00681f
C2277 avdd.n1233 dvss 0.460184f
C2278 avdd.n1235 dvss 0.286865f
C2279 avdd.n1237 dvss 0.286865f
C2280 avdd.n1239 dvss 0.326308f
C2281 avdd.n1241 dvss 0.326308f
C2282 avdd.n1243 dvss 0.286865f
C2283 avdd.n1245 dvss 0.286865f
C2284 avdd.n1247 dvss 0.286865f
C2285 avdd.n1249 dvss 0.286865f
C2286 avdd.n1251 dvss 0.286865f
C2287 avdd.n1253 dvss 0.258624f
C2288 avdd.n1254 dvss 0.115125f
C2289 avdd.n1256 dvss 0.247668f
C2290 avdd.n1257 dvss 2.57803f
C2291 avdd.n1258 dvss 0.880834f
C2292 avdd.n1259 dvss 0.978922f
C2293 avdd.n1260 dvss 0.993149f
C2294 avdd.n1261 dvss 4.22301f
C2295 avdd.n1262 dvss 4.22247f
C2296 avdd.n1263 dvss 15.931701f
C2297 avdd.n1264 dvss 1.02641f
C2298 avdd.n1265 dvss 0.99239f
C2299 avdd.n1266 dvss 0.901373f
C2300 avdd.n1267 dvss 1.80268f
C2301 avdd.n1268 dvss 0.880834f
C2302 avdd.n1269 dvss 1.53938f
C2303 avdd.n1270 dvss 0.115125f
C2304 avdd.n1271 dvss 0.142138f
C2305 avdd.n1272 dvss 0.136266f
C2306 avdd.n1273 dvss 0.127835f
C2307 avdd.n1274 dvss 0.78481f
C2308 avdd.n1275 dvss 2.8425f
C2309 avdd.n1276 dvss 3.13648f
C2310 avdd.n1277 dvss 2.83597f
C2311 avdd.n1278 dvss 0.794727f
C2312 avdd.n1279 dvss 0.166768f
C2313 avdd.n1280 dvss 0.236203f
C2314 avdd.t590 dvss 0.704956f
C2315 avdd.n1281 dvss 0.539054f
C2316 avdd.t598 dvss 0.704956f
C2317 avdd.t586 dvss 0.939941f
C2318 avdd.t600 dvss 0.939941f
C2319 avdd.t596 dvss 0.939941f
C2320 avdd.t592 dvss 1.1627f
C2321 avdd.n1282 dvss 1.5397f
C2322 avdd.t588 dvss 0.939941f
C2323 avdd.t594 dvss 0.939941f
C2324 avdd.t604 dvss 0.939941f
C2325 avdd.t602 dvss 1.1627f
C2326 avdd.n1283 dvss 1.5397f
C2327 avdd.n1284 dvss 0.18791f
C2328 avdd.n1285 dvss 0.172686f
C2329 avdd.n1286 dvss 0.317697f
C2330 avdd.n1287 dvss 0.172686f
C2331 avdd.n1289 dvss 0.286865f
C2332 avdd.n1291 dvss 0.286865f
C2333 avdd.n1293 dvss 0.286865f
C2334 avdd.n1295 dvss 0.286865f
C2335 avdd.n1297 dvss 0.286865f
C2336 avdd.n1299 dvss 0.326308f
C2337 avdd.n1301 dvss 0.326308f
C2338 avdd.n1303 dvss 0.286865f
C2339 avdd.n1305 dvss 0.286865f
C2340 avdd.n1307 dvss 0.460184f
C2341 avdd.n1308 dvss 3.62023f
C2342 avdd.n1309 dvss 2.72536f
C2343 avdd.n1310 dvss 0.170379f
C2344 avdd.n1311 dvss 0.326308f
C2345 avdd.t354 dvss 2.85263f
C2346 avdd.n1312 dvss 0.170379f
C2347 avdd.n1313 dvss 0.286865f
C2348 avdd.t271 dvss 2.85333f
C2349 avdd.n1314 dvss 0.170379f
C2350 avdd.t269 dvss 2.85333f
C2351 avdd.n1315 dvss 1.40632f
C2352 avdd.n1317 dvss 0.258624f
C2353 avdd.t300 dvss 2.85333f
C2354 avdd.n1318 dvss 1.40632f
C2355 avdd.n1320 dvss 0.286865f
C2356 avdd.n1321 dvss 0.286865f
C2357 avdd.t307 dvss 2.85333f
C2358 avdd.n1323 dvss 1.40632f
C2359 avdd.n1324 dvss 0.170379f
C2360 avdd.t325 dvss 2.85333f
C2361 avdd.n1326 dvss 1.40632f
C2362 avdd.n1327 dvss 0.170379f
C2363 avdd.n1328 dvss 0.170379f
C2364 avdd.n1329 dvss 1.40632f
C2365 avdd.n1331 dvss 0.286865f
C2366 avdd.t330 dvss 2.85333f
C2367 avdd.n1332 dvss 1.40632f
C2368 avdd.n1334 dvss 0.286865f
C2369 avdd.n1335 dvss 0.326308f
C2370 avdd.t275 dvss 2.85333f
C2371 avdd.n1337 dvss 1.40632f
C2372 avdd.n1338 dvss 0.209822f
C2373 avdd.t346 dvss 2.85263f
C2374 avdd.n1340 dvss 1.4013f
C2375 avdd.n1341 dvss 0.209822f
C2376 avdd.n1342 dvss 0.170379f
C2377 avdd.n1343 dvss 1.4013f
C2378 avdd.n1345 dvss 0.286865f
C2379 avdd.t348 dvss 2.85263f
C2380 avdd.n1346 dvss 1.4013f
C2381 avdd.n1348 dvss 0.286865f
C2382 avdd.n1349 dvss 0.460184f
C2383 avdd.t364 dvss 2.85263f
C2384 avdd.n1351 dvss 1.4013f
C2385 avdd.n1352 dvss 0.343698f
C2386 avdd.n1353 dvss 2.01084f
C2387 avdd.n1354 dvss 0.830753f
C2388 avdd.n1355 dvss 0.241516f
C2389 avdd.n1357 dvss 0.285283f
C2390 avdd.n1359 dvss 0.285283f
C2391 avdd.n1361 dvss 0.285283f
C2392 avdd.n1363 dvss 0.285283f
C2393 avdd.n1364 dvss 0.306627f
C2394 avdd.n1365 dvss 0.189145f
C2395 avdd.n1366 dvss 0.289183f
C2396 avdd.n1367 dvss 0.539054f
C2397 avdd.n1368 dvss 2.22853f
C2398 avdd.n1369 dvss 0.563898f
C2399 avdd.t140 dvss 61.383f
C2400 avdd.t240 dvss 48.5178f
C2401 avdd.n1370 dvss 0.834636f
C2402 avdd.n1371 dvss 1.42313f
C2403 avdd.n1372 dvss 19.5848f
C2404 avdd.n1373 dvss 1.19282f
C2405 avdd.n1374 dvss 0.713752f
C2406 avdd.n1375 dvss 0.217503f
C2407 avdd.n1376 dvss 0.247032f
C2408 avdd.n1377 dvss 0.115125f
C2409 avdd.n1378 dvss 0.213134f
C2410 avdd.t239 dvss 2.86945f
C2411 avdd.n1379 dvss 1.3892f
C2412 avdd.n1381 dvss 0.794824f
C2413 avdd.n1382 dvss 2.04908f
C2414 avdd.n1383 dvss 2.50608f
C2415 avdd.n1384 dvss 1.96847f
C2416 avdd.n1385 dvss 0.960954f
C2417 avdd.n1386 dvss 0.980125f
C2418 avdd.n1387 dvss 4.23964f
C2419 avdd.n1388 dvss 16.1996f
C2420 avdd.n1389 dvss 15.9296f
C2421 avdd.n1390 dvss 16.1996f
C2422 avdd.n1391 dvss 4.23964f
C2423 avdd.n1392 dvss 0.979544f
C2424 avdd.n1393 dvss 0.948763f
C2425 avdd.n1394 dvss 1.96847f
C2426 avdd.n1395 dvss 1.77298f
C2427 avdd.n1396 dvss 1.95878f
C2428 avdd.n1397 dvss 0.637456f
C2429 avdd.n1398 dvss 1.16091f
C2430 avdd.n1399 dvss 1.93485f
C2431 avdd.n1400 dvss 0.605048f
C2432 avdd.n1402 dvss 0.2402f
C2433 avdd.n1403 dvss 0.115125f
C2434 avdd.n1404 dvss 0.846056f
C2435 avdd.n1405 dvss 2.16083f
C2436 avdd.n1406 dvss 30.6915f
C2437 avdd.n1407 dvss 2.16083f
C2438 avdd.n1408 dvss 1.26669f
C2439 avdd.n1409 dvss 0.771102f
C2440 avdd.n1410 dvss 0.834636f
C2441 avdd.n1411 dvss 1.42313f
C2442 avdd.n1412 dvss 19.5848f
C2443 avdd.n1413 dvss 1.19282f
C2444 avdd.n1414 dvss 0.713752f
C2445 avdd.n1415 dvss 0.14348f
C2446 avdd.n1416 dvss 0.247032f
C2447 avdd.n1417 dvss 0.115125f
C2448 avdd.t304 dvss 2.85333f
C2449 avdd.n1418 dvss 1.40632f
C2450 avdd.n1419 dvss 0.142138f
C2451 avdd.t356 dvss 2.85333f
C2452 avdd.n1420 dvss 1.40632f
C2453 avdd.n1421 dvss 0.170379f
C2454 avdd.t359 dvss 2.85333f
C2455 avdd.n1422 dvss 1.40632f
C2456 avdd.n1423 dvss 0.170379f
C2457 avdd.t377 dvss 2.85333f
C2458 avdd.n1424 dvss 1.40632f
C2459 avdd.n1425 dvss 0.170379f
C2460 avdd.t235 dvss 2.85333f
C2461 avdd.n1426 dvss 1.40632f
C2462 avdd.n1427 dvss 0.170379f
C2463 avdd.t284 dvss 2.85333f
C2464 avdd.n1428 dvss 1.40632f
C2465 avdd.n1429 dvss 0.170379f
C2466 avdd.t242 dvss 2.85333f
C2467 avdd.n1430 dvss 1.40632f
C2468 avdd.n1431 dvss 0.209822f
C2469 avdd.t291 dvss 2.85263f
C2470 avdd.n1432 dvss 1.4013f
C2471 avdd.n1433 dvss 0.209822f
C2472 avdd.t311 dvss 2.85263f
C2473 avdd.n1434 dvss 1.4013f
C2474 avdd.n1435 dvss 0.170379f
C2475 avdd.t297 dvss 2.85263f
C2476 avdd.n1436 dvss 1.4013f
C2477 avdd.n1437 dvss 0.170379f
C2478 avdd.t320 dvss 2.85263f
C2479 avdd.n1438 dvss 1.4013f
C2480 avdd.n1439 dvss 0.343698f
C2481 avdd.n1440 dvss 1.32207f
C2482 avdd.n1441 dvss 0.516245f
C2483 avdd.n1442 dvss 1.04548f
C2484 avdd.n1443 dvss 0.774177f
C2485 avdd.n1444 dvss 3.19868f
C2486 avdd.n1445 dvss 5.19383f
C2487 avdd.n1446 dvss 2.97397f
C2488 avdd.n1447 dvss 1.92291f
C2489 avdd.n1448 dvss 13.0557f
C2490 avdd.n1449 dvss 9.19242f
C2491 avdd.n1450 dvss 50.164803f
C2492 avdd.n1451 dvss 42.835197f
C2493 avdd.n1452 dvss 4.38592f
C2494 avdd.n1453 dvss 4.69133f
C2495 avdd.n1454 dvss 1.06368f
C2496 avdd.n1455 dvss 6.50313f
C2497 avdd.n1456 dvss 2.29325f
C2498 avdd.n1457 dvss 8.80394f
C2499 avdd.n1458 dvss 14.4214f
C2500 avdd.n1459 dvss 3.70579f
C2501 avdd.n1460 dvss 0.655638f
C2502 avdd.n1461 dvss 1.75246f
C2503 avdd.n1462 dvss 7.12364f
C2504 avdd.n1463 dvss 1.42958f
C2505 avdd.n1464 dvss 7.95466f
C2506 avdd.n1465 dvss 2.22993f
C2507 avdd.n1466 dvss 2.23103f
C2508 avdd.n1467 dvss 27.336699f
C2509 avdd.n1468 dvss 7.13531f
C2510 avdd.n1469 dvss 1.0444f
C2511 avdd.n1470 dvss 1.04895f
C2512 avdd.n1471 dvss 3.72287f
C2513 avdd.n1472 dvss 3.68745f
C2514 avdd.n1473 dvss 1.75636f
C2515 avdd.n1474 dvss 0.65743f
C2516 avdd.n1475 dvss 5.25296f
C2517 avdd.n1476 dvss 20.6425f
C2518 avdd.n1477 dvss 33.9332f
C2519 avdd.n1478 dvss 41.8823f
C2520 avdd.n1479 dvss 10.113299f
C2521 avdd.n1480 dvss 2.29244f
C2522 avdd.n1481 dvss 2.66377f
C2523 avdd.n1482 dvss 10.7805f
C2524 avdd.n1483 dvss 10.0564f
C2525 avdd.n1484 dvss 5.29402f
C2526 avdd.n1485 dvss 2.43554f
C2527 avdd.n1486 dvss 1.61378f
C2528 avdd.n1487 dvss 5.82401f
C2529 avdd.n1488 dvss 6.72044f
C2530 avdd.n1489 dvss 1.06674f
C2531 avdd.n1490 dvss 2.03649f
C2532 avdd.n1491 dvss 5.25803f
C2533 avdd.n1492 dvss 27.169802f
C2534 avdd.n1493 dvss 35.232998f
C2535 avdd.n1494 dvss 57.8455f
C2536 avdd.n1495 dvss 15.063001f
C2537 avdd.n1496 dvss 1.49167f
C2538 avdd.n1497 dvss 2.33649f
C2539 avdd.n1498 dvss 6.49862f
C2540 avdd.n1499 dvss 3.75552f
C2541 avdd.n1500 dvss 30.6886f
C2542 avdd.n1501 dvss 71.7888f
C2543 avdd.n1502 dvss 8.9529f
C2544 avdd.n1503 dvss 1.94835f
C2545 avdd.t345 dvss 0.105757f
C2546 avdd.t572 dvss 0.105757f
C2547 avdd.n1504 dvss 0.268539f
C2548 avdd.n1505 dvss 0.599458f
C2549 avdd.n1506 dvss 1.48879f
C2550 avdd.n1507 dvss 1.39103f
C2551 avdd.n1508 dvss 0.218054f
C2552 avdd.n1509 dvss 0.290937f
C2553 avdd.n1510 dvss 0.610642f
C2554 avdd.n1511 dvss 0.694497f
C2555 avdd.t217 dvss 4.63479f
C2556 avdd.t448 dvss 2.3174f
C2557 avdd.n1512 dvss 0.610642f
C2558 avdd.n1514 dvss 0.308118f
C2559 avdd.n1515 dvss 0.523075f
C2560 avdd.t100 dvss 5.96274f
C2561 avdd.t234 dvss 4.63479f
C2562 avdd.t220 dvss 4.63479f
C2563 avdd.t163 dvss 3.12458f
C2564 avdd.t446 dvss 2.90326f
C2565 avdd.n1516 dvss 0.284699f
C2566 avdd.n1517 dvss 6.822f
C2567 avdd.t569 dvss 9.0743f
C2568 avdd.t96 dvss 5.96274f
C2569 avdd.t555 dvss 7.577109f
C2570 avdd.n1518 dvss 0.523075f
C2571 avdd.n1519 dvss 1.53444f
C2572 avdd.t575 dvss 0.443137f
C2573 avdd.n1520 dvss 1.09699f
C2574 avdd.t548 dvss 0.443137f
C2575 avdd.n1521 dvss 0.956185f
C2576 avdd.t343 dvss 0.885595f
C2577 avdd.n1522 dvss 0.802714f
C2578 avdd.t350 dvss 0.88547f
C2579 avdd.n1523 dvss 0.950446f
C2580 avdd.t233 dvss 0.88547f
C2581 avdd.n1524 dvss 1.06973f
C2582 avdd.n1525 dvss 0.163797f
C2583 avdd.n1526 dvss 0.496155f
C2584 avdd.t570 dvss 0.443137f
C2585 avdd.n1527 dvss 1.03391f
C2586 avdd.t546 dvss 0.105757f
C2587 avdd.t556 dvss 0.105757f
C2588 avdd.n1528 dvss 0.270278f
C2589 avdd.n1529 dvss 1.41624f
C2590 avdd.t558 dvss 0.105757f
C2591 avdd.t219 dvss 0.105757f
C2592 avdd.n1530 dvss 0.270278f
C2593 avdd.n1531 dvss 1.24137f
C2594 avdd.n1532 dvss 0.503171f
C2595 avdd.n1533 dvss 0.163797f
C2596 avdd.n1534 dvss 0.293649f
C2597 avdd.t323 dvss 1.43218f
C2598 avdd.n1535 dvss 2.98705f
C2599 avdd.t574 dvss 3.19062f
C2600 avdd.t218 dvss 8.33221f
C2601 avdd.t557 dvss 8.8009f
C2602 avdd.t231 dvss 4.72593f
C2603 avdd.n1537 dvss 0.284699f
C2604 avdd.n1538 dvss 5.31179f
C2605 avdd.t547 dvss 5.44198f
C2606 avdd.n1539 dvss 3.24721f
C2607 avdd.n1540 dvss 3.24721f
C2608 avdd.n1541 dvss 1.90495f
C2609 avdd.n1542 dvss 1.88493f
C2610 avdd.n1543 dvss 1.8255f
C2611 avdd.t573 dvss 3.54119f
C2612 avdd.t344 dvss 4.63479f
C2613 avdd.t571 dvss 4.63479f
C2614 avdd.t164 dvss 5.22065f
C2615 avdd.n1544 dvss 2.99439f
C2616 avdd.t94 dvss 6.64951f
C2617 avdd.t90 dvss 9.67256f
C2618 avdd.t92 dvss 7.48133f
C2619 avdd.n1545 dvss 4.98756f
C2620 avdd.t98 dvss 7.48133f
C2621 avdd.t336 dvss 9.975111f
C2622 avdd.t505 dvss 9.975111f
C2623 avdd.t507 dvss 9.975111f
C2624 avdd.t371 dvss 9.975111f
C2625 avdd.t509 dvss 9.975111f
C2626 avdd.t511 dvss 9.975111f
C2627 avdd.t264 dvss 8.39037f
C2628 avdd.n1546 dvss 7.51454f
C2629 avdd.n1547 dvss 0.971795f
C2630 avdd.n1548 dvss 0.980201f
C2631 avdd.n1549 dvss 2.95326f
C2632 avdd.t335 dvss 4.46957f
C2633 avdd.n1550 dvss 1.65121f
C2634 avdd.n1551 dvss 1.82683f
C2635 avdd.n1552 dvss 0.364135f
C2636 avdd.t266 dvss 0.391979f
C2637 avdd.t263 dvss 4.57993f
C2638 avdd.n1553 dvss 4.05933f
C2639 avdd.n1554 dvss 0.728002f
C2640 avdd.t512 dvss 0.105757f
C2641 avdd.t265 dvss 0.105757f
C2642 avdd.n1555 dvss 0.225995f
C2643 avdd.n1556 dvss 1.49865f
C2644 avdd.n1557 dvss 1.49865f
C2645 avdd.t508 dvss 0.105757f
C2646 avdd.t510 dvss 0.105757f
C2647 avdd.n1558 dvss 0.225995f
C2648 avdd.t372 dvss 0.211515f
C2649 avdd.n1559 dvss 0.217774f
C2650 avdd.t370 dvss 4.57171f
C2651 avdd.n1560 dvss 4.03021f
C2652 avdd.n1561 dvss 1.43681f
C2653 avdd.t99 dvss 0.105757f
C2654 avdd.n1562 dvss 0.215426f
C2655 avdd.t337 dvss 0.211515f
C2656 avdd.t506 dvss 0.105757f
C2657 avdd.n1563 dvss 0.225995f
C2658 avdd.n1564 dvss 1.49919f
C2659 avdd.n1565 dvss 1.03187f
C2660 avdd.n1566 dvss 0.171066f
C2661 avdd.n1567 dvss 1.81475f
C2662 avdd.n1568 dvss 1.62776f
C2663 avdd.n1569 dvss 1.80208f
C2664 avdd.t91 dvss 0.105757f
C2665 avdd.t93 dvss 0.105757f
C2666 avdd.n1570 dvss 0.225995f
C2667 avdd.n1571 dvss 1.42525f
C2668 avdd.t449 dvss 0.105757f
C2669 avdd.t95 dvss 0.105757f
C2670 avdd.n1572 dvss 0.225995f
C2671 avdd.n1573 dvss 1.96174f
C2672 avdd.t97 dvss 0.105757f
C2673 avdd.t447 dvss 0.105757f
C2674 avdd.n1574 dvss 0.225995f
C2675 avdd.n1575 dvss 1.96174f
C2676 avdd.n1576 dvss 1.49865f
C2677 avdd.t101 dvss 0.105757f
C2678 avdd.n1577 dvss 0.225995f
C2679 avdd.t232 dvss 0.497736f
C2680 avdd.t230 dvss 4.57993f
C2681 avdd.n1578 dvss 4.05933f
C2682 avdd.n1579 dvss 0.724799f
C2683 avdd.n1580 dvss 3.3406f
C2684 avdd.n1581 dvss 0.980201f
C2685 avdd.n1582 dvss 0.971795f
C2686 avdd.n1583 dvss 3.26744f
C2687 avdd.n1584 dvss 3.3311f
C2688 avdd.n1585 dvss 0.216527f
C2689 avdd.n1586 dvss 0.369662f
C2690 avdd.t324 dvss 2.75325f
C2691 avdd.n1587 dvss 0.369662f
C2692 avdd.n1588 dvss 0.664432f
C2693 avdd.n1589 dvss 0.283692f
C2694 avdd.n1590 dvss 0.158585f
C2695 avdd.n1591 dvss 0.209917f
C2696 avdd.n1592 dvss 0.541054f
C2697 avdd.t545 dvss 9.556009f
C2698 avdd.n1593 dvss 0.541054f
C2699 avdd.n1594 dvss 0.209917f
C2700 avdd.n1595 dvss 0.158585f
C2701 avdd.n1596 dvss 0.308118f
C2702 avdd.n1597 dvss 0.31858f
C2703 avdd.n1598 dvss 0.543016f
C2704 avdd.t351 dvss 3.411f
C2705 avdd.n1599 dvss 0.543016f
C2706 avdd.n1600 dvss 0.300735f
C2707 avdd.n1601 dvss 0.234397f
C2708 avdd.n1602 dvss 1.53339f
C2709 avdd.n1603 dvss 2.22509f
C2710 avdd.n1604 dvss 14.7798f
C2711 avdd.n1605 dvss 31.0439f
C2712 avdd.n1606 dvss 20.1994f
C2713 avdd.t59 dvss 0.469755f
C2714 avdd.n1607 dvss 0.89587f
C2715 avdd.n1608 dvss 0.772198f
C2716 avdd.n1609 dvss 0.311548f
C2717 avdd.t73 dvss 0.105757f
C2718 avdd.t89 dvss 0.105757f
C2719 avdd.n1610 dvss 0.299286f
C2720 avdd.n1611 dvss 0.974644f
C2721 avdd.t69 dvss 0.105757f
C2722 avdd.t85 dvss 0.105757f
C2723 avdd.n1612 dvss 0.299286f
C2724 avdd.n1613 dvss 0.974644f
C2725 avdd.t81 dvss 0.105757f
C2726 avdd.t63 dvss 0.105757f
C2727 avdd.n1614 dvss 0.299286f
C2728 avdd.n1615 dvss 0.974644f
C2729 avdd.t77 dvss 0.105757f
C2730 avdd.t61 dvss 0.105757f
C2731 avdd.n1616 dvss 0.299286f
C2732 avdd.n1617 dvss 0.974644f
C2733 avdd.t75 dvss 0.105757f
C2734 avdd.t71 dvss 0.105757f
C2735 avdd.n1618 dvss 0.299286f
C2736 avdd.n1619 dvss 0.974644f
C2737 avdd.t87 dvss 0.105757f
C2738 avdd.t67 dvss 0.105757f
C2739 avdd.n1620 dvss 0.299286f
C2740 avdd.n1621 dvss 0.974644f
C2741 avdd.t83 dvss 0.105757f
C2742 avdd.t65 dvss 0.105757f
C2743 avdd.n1622 dvss 0.299286f
C2744 avdd.n1623 dvss 0.974644f
C2745 avdd.t79 dvss 0.469755f
C2746 avdd.n1624 dvss 1.03881f
C2747 avdd.n1625 dvss 1.01983f
C2748 avdd.n1626 dvss 0.319252f
C2749 avdd.n1627 dvss 0.9361f
C2750 avdd.n1628 dvss 0.311548f
C2751 avdd.n1629 dvss 0.451432f
C2752 avdd.n1630 dvss 0.9361f
C2753 avdd.n1631 dvss 3.07507f
C2754 avdd.t58 dvss 2.39529f
C2755 avdd.t72 dvss 1.97855f
C2756 avdd.t88 dvss 1.97855f
C2757 avdd.t68 dvss 1.97855f
C2758 avdd.t84 dvss 1.97855f
C2759 avdd.t80 dvss 1.97855f
C2760 avdd.t62 dvss 1.97855f
C2761 avdd.t76 dvss 1.48391f
C2762 avdd.n1632 dvss 0.989275f
C2763 avdd.t60 dvss 1.48391f
C2764 avdd.t74 dvss 1.97855f
C2765 avdd.t70 dvss 1.97855f
C2766 avdd.t86 dvss 1.97855f
C2767 avdd.t66 dvss 1.97855f
C2768 avdd.t82 dvss 1.97855f
C2769 avdd.t64 dvss 1.97855f
C2770 avdd.t78 dvss 2.39529f
C2771 avdd.n1633 dvss 3.07507f
C2772 avdd.n1634 dvss 0.319252f
C2773 avdd.n1635 dvss 0.550028f
C2774 avdd.n1636 dvss 1.08605f
C2775 avdd.n1637 dvss 1.01875f
C2776 avdd.n1638 dvss 0.370514f
C2777 avdd.n1639 dvss 1.38238f
C2778 avdd.n1640 dvss 1.16827f
C2779 avdd.n1641 dvss 1.0953f
C2780 avdd.n1642 dvss 1.8195f
C2781 avdd.n1643 dvss 1.09168f
C2782 avdd.n1644 dvss 0.63618f
C2783 avdd.n1645 dvss 0.15869f
C2784 avdd.n1646 dvss 4.24618f
C2785 avdd.t492 dvss 2.39529f
C2786 avdd.t491 dvss 1.97855f
C2787 avdd.t310 dvss 1.97855f
C2788 avdd.t156 dvss 1.97855f
C2789 avdd.t155 dvss 1.97855f
C2790 avdd.t249 dvss 1.97855f
C2791 avdd.t180 dvss 1.97855f
C2792 avdd.t179 dvss 1.97855f
C2793 avdd.t339 dvss 1.97855f
C2794 avdd.t504 dvss 1.97855f
C2795 avdd.t503 dvss 1.97855f
C2796 avdd.t281 dvss 1.97855f
C2797 avdd.t522 dvss 1.97855f
C2798 avdd.t523 dvss 1.97855f
C2799 avdd.t381 dvss 1.97855f
C2800 avdd.t109 dvss 1.97855f
C2801 avdd.t108 dvss 1.97855f
C2802 avdd.t268 dvss 1.97855f
C2803 avdd.t152 dvss 1.97855f
C2804 avdd.t151 dvss 1.97855f
C2805 avdd.t399 dvss 1.97855f
C2806 avdd.t420 dvss 1.97855f
C2807 avdd.t419 dvss 1.97855f
C2808 avdd.t387 dvss 1.97855f
C2809 avdd.t170 dvss 1.97855f
C2810 avdd.t171 dvss 1.97855f
C2811 avdd.t374 dvss 1.97855f
C2812 avdd.t490 dvss 1.97855f
C2813 avdd.t489 dvss 1.97855f
C2814 avdd.t385 dvss 1.97855f
C2815 avdd.t167 dvss 1.97855f
C2816 avdd.t168 dvss 1.97855f
C2817 avdd.t303 dvss 1.97855f
C2818 avdd.t402 dvss 1.97855f
C2819 avdd.t403 dvss 1.97855f
C2820 avdd.t397 dvss 1.97855f
C2821 avdd.t499 dvss 1.97855f
C2822 avdd.t500 dvss 1.97855f
C2823 avdd.t401 dvss 1.97855f
C2824 avdd.t2 dvss 1.97855f
C2825 avdd.t3 dvss 1.97855f
C2826 avdd.t363 dvss 1.97855f
C2827 avdd.t214 dvss 1.97855f
C2828 avdd.t213 dvss 1.97855f
C2829 avdd.t254 dvss 1.97855f
C2830 avdd.t412 dvss 1.97855f
C2831 avdd.t413 dvss 2.39529f
C2832 avdd.n1647 dvss 4.24618f
C2833 avdd.n1648 dvss 0.158982f
C2834 avdd.n1649 dvss 0.635391f
C2835 avdd.n1650 dvss 0.297765f
C2836 avdd.n1651 dvss 1.3008f
C2837 avdd.n1652 dvss 0.989319f
C2838 rstring_mux_0.vtrip4.t9 dvss 0.171176f
C2839 rstring_mux_0.vtrip4.n0 dvss 0.18541f
C2840 rstring_mux_0.vtrip4.n1 dvss 0.121565f
C2841 rstring_mux_0.vtrip4.n2 dvss 1.18871f
C2842 rstring_mux_0.vtrip4.n3 dvss 0.18541f
C2843 rstring_mux_0.vtrip4.n4 dvss 0.121565f
C2844 rstring_mux_0.vtrip4.n5 dvss 0.749847f
C2845 rstring_mux_0.vtrip4.n6 dvss 1.88677f
C2846 rstring_mux_0.vtrip4.n7 dvss 2.28683f
C2847 rstring_mux_0.vtrip4.t0 dvss 0.726836f
C2848 vin_vunder.n0 dvss 0.115783f
C2849 vin_vunder.n1 dvss 0.128888f
C2850 vin_vunder.n2 dvss 0.116135f
C2851 vin_vunder.n3 dvss 0.316141f
C2852 vin_vunder.n4 dvss 0.316141f
C2853 vin_vunder.n5 dvss 0.316141f
C2854 vin_vunder.n6 dvss 0.128888f
C2855 vin_vunder.n7 dvss 0.272716f
C2856 vin_vunder.n8 dvss 0.116135f
C2857 vin_vunder.n9 dvss 0.128888f
C2858 vin_vunder.n10 dvss 0.27262f
C2859 vin_vunder.n11 dvss 0.12947f
C2860 vin_vunder.n12 dvss 0.116135f
C2861 vin_vunder.n13 dvss 0.128888f
C2862 vin_vunder.n14 dvss 0.27262f
C2863 vin_vunder.n15 dvss 0.131247f
C2864 vin_vunder.n16 dvss -0.538117f
C2865 vin_vunder.n17 dvss 0.624066f
C2866 vin_vunder.n18 dvss 0.12947f
C2867 vin_vunder.n19 dvss 0.27262f
C2868 vin_vunder.n20 dvss 0.128888f
C2869 vin_vunder.n21 dvss 0.116135f
C2870 vin_vunder.n22 dvss 0.316141f
C2871 vin_vunder.n23 dvss 0.157318f
C2872 vin_vunder.t56 dvss 2.07495f
C2873 vin_vunder.t53 dvss 1.98572f
C2874 vin_vunder.n24 dvss 1.65357f
C2875 vin_vunder.t61 dvss 1.98572f
C2876 vin_vunder.n25 dvss 0.873349f
C2877 vin_vunder.t58 dvss 1.98572f
C2878 vin_vunder.n26 dvss 0.873349f
C2879 vin_vunder.t49 dvss 1.98572f
C2880 vin_vunder.n27 dvss 0.873349f
C2881 vin_vunder.t59 dvss 1.98572f
C2882 vin_vunder.n28 dvss 0.873349f
C2883 vin_vunder.t55 dvss 1.98572f
C2884 vin_vunder.n29 dvss 0.873349f
C2885 vin_vunder.t54 dvss 1.98572f
C2886 vin_vunder.n30 dvss 1.03295f
C2887 vin_vunder.t50 dvss 2.0927f
C2888 vin_vunder.t62 dvss 2.00221f
C2889 vin_vunder.n31 dvss 1.69074f
C2890 vin_vunder.t57 dvss 2.00221f
C2891 vin_vunder.n32 dvss 0.892563f
C2892 vin_vunder.t51 dvss 2.00221f
C2893 vin_vunder.n33 dvss 0.892563f
C2894 vin_vunder.t60 dvss 2.00221f
C2895 vin_vunder.n34 dvss 0.892563f
C2896 vin_vunder.t52 dvss 2.00221f
C2897 vin_vunder.n35 dvss 0.892563f
C2898 vin_vunder.t48 dvss 2.00221f
C2899 vin_vunder.n36 dvss 0.892563f
C2900 vin_vunder.t63 dvss 2.00221f
C2901 vin_vunder.n37 dvss 0.987086f
C2902 vin_vunder.n38 dvss 3.5161f
C2903 vin_vunder.n39 dvss 3.47781f
C2904 vin_vunder.n40 dvss 0.291279f
C2905 vin_vunder.n41 dvss 0.147063f
C2906 vin_vunder.n42 dvss 0.158436f
C2907 vin_vunder.n43 dvss 0.572763f
C2908 vin_vunder.n44 dvss 0.147063f
C2909 vin_vunder.n45 dvss 0.158436f
C2910 vin_vunder.n46 dvss 0.572763f
C2911 vin_vunder.n47 dvss 0.147063f
C2912 vin_vunder.n48 dvss 0.158436f
C2913 vin_vunder.n49 dvss 0.572763f
C2914 vin_vunder.n50 dvss 0.147063f
C2915 vin_vunder.n51 dvss 0.158436f
C2916 vin_vunder.n52 dvss 0.572763f
C2917 vin_vunder.n53 dvss 0.316141f
C2918 vin_vunder.n54 dvss 0.281145f
C2919 vin_vunder.n55 dvss 0.116135f
C2920 vin_vunder.n56 dvss 0.128888f
C2921 vin_vunder.n57 dvss 0.147063f
C2922 vin_vunder.n58 dvss 0.158436f
C2923 vin_vunder.n59 dvss 0.572763f
C2924 vin_vunder.n60 dvss 0.147063f
C2925 vin_vunder.n61 dvss 0.158436f
C2926 vin_vunder.t29 dvss 0.196899f
C2927 vin_vunder.n62 dvss 0.334106f
C2928 vin_vunder.t44 dvss 0.213769f
C2929 vin_vunder.n63 dvss 0.604784f
C2930 vin_vunder.n64 dvss 0.158436f
C2931 vin_vunder.n65 dvss 0.147063f
C2932 vin_vunder.n66 dvss 0.572763f
C2933 vin_vunder.n67 dvss 0.128888f
C2934 vin_vunder.n68 dvss 0.116135f
C2935 vin_vunder.n69 dvss 0.316141f
C2936 vin_vunder.n70 dvss 0.27262f
C2937 vin_vunder.n71 dvss 0.206988f
C2938 vin_vunder.n72 dvss 0.12947f
C2939 vin_vunder.n73 dvss 0.27262f
C2940 vin_vunder.n74 dvss 0.128888f
C2941 vin_vunder.n75 dvss 0.116135f
C2942 vin_vunder.n76 dvss 0.316141f
C2943 vin_vunder.n77 dvss 0.27262f
C2944 avss.n1 dvss 0.652329f
C2945 avss.n7 dvss 2.70631f
C2946 avss.t254 dvss 7.02941f
C2947 avss.n8 dvss 13.955701f
C2948 avss.t204 dvss 6.73382f
C2949 avss.n9 dvss 0.210222f
C2950 avss.n10 dvss 0.210222f
C2951 avss.n11 dvss 0.295554f
C2952 avss.t88 dvss 0.464418f
C2953 avss.t186 dvss 6.73382f
C2954 avss.t252 dvss 9.2942f
C2955 avss.n12 dvss 0.299831f
C2956 avss.n13 dvss 0.299831f
C2957 avss.n14 dvss 0.176051f
C2958 avss.n15 dvss 0.146585f
C2959 avss.t316 dvss 0.221192f
C2960 avss.t299 dvss 0.216631f
C2961 avss.n16 dvss 0.882838f
C2962 avss.n17 dvss 0.208683f
C2963 avss.t317 dvss 9.67826f
C2964 avss.t201 dvss 11.7266f
C2965 avss.t165 dvss 9.67826f
C2966 avss.t158 dvss 5.86329f
C2967 avss.n18 dvss 9.67826f
C2968 avss.t326 dvss 5.86329f
C2969 avss.t163 dvss 9.67826f
C2970 avss.t179 dvss 9.65266f
C2971 avss.t141 dvss 3.53333f
C2972 avss.t196 dvss 8.21884f
C2973 avss.t151 dvss 9.2942f
C2974 avss.t304 dvss 5.58164f
C2975 avss.n19 dvss 0.401911f
C2976 avss.n20 dvss 0.401911f
C2977 avss.n21 dvss 0.236133f
C2978 avss.n22 dvss 0.131025f
C2979 avss.t53 dvss 0.355198f
C2980 avss.n23 dvss 0.348225f
C2981 avss.t81 dvss 0.355217f
C2982 avss.n24 dvss 0.301805f
C2983 avss.t9 dvss 0.355201f
C2984 avss.n25 dvss 0.657754f
C2985 avss.n26 dvss 2.06181f
C2986 avss.n27 dvss 1.04504f
C2987 avss.t15 dvss 4.16156f
C2988 avss.t18 dvss 0.16157f
C2989 avss.n28 dvss 1.57106f
C2990 avss.n29 dvss 0.407738f
C2991 avss.n30 dvss 0.650677f
C2992 avss.n31 dvss 0.153488f
C2993 avss.n32 dvss 0.165885f
C2994 avss.n33 dvss 1.27521f
C2995 avss.n34 dvss 1.27521f
C2996 avss.t37 dvss 4.16156f
C2997 avss.n35 dvss 0.165885f
C2998 avss.t38 dvss 0.204737f
C2999 avss.n36 dvss 1.57106f
C3000 avss.n37 dvss 0.466083f
C3001 avss.n38 dvss 0.459112f
C3002 avss.n40 dvss 0.938505f
C3003 avss.t48 dvss 4.16156f
C3004 avss.t50 dvss 0.16157f
C3005 avss.n41 dvss 1.57106f
C3006 avss.n42 dvss 0.407738f
C3007 avss.n44 dvss 0.703565f
C3008 avss.n45 dvss 0.703565f
C3009 avss.t315 dvss 2.09951f
C3010 avss.t298 dvss 9.67826f
C3011 avss.t199 dvss 6.6058f
C3012 avss.t89 dvss 7.57874f
C3013 avss.n46 dvss 6.6058f
C3014 avss.n47 dvss 1.10961f
C3015 avss.n48 dvss 1.10961f
C3016 avss.n49 dvss 8.42142f
C3017 avss.t198 dvss 4.94155f
C3018 avss.n50 dvss 1.75259f
C3019 avss.n51 dvss 1.75259f
C3020 avss.n52 dvss 1.75259f
C3021 avss.n53 dvss 2.78345f
C3022 avss.n54 dvss 1.75444f
C3023 avss.n55 dvss 0.14706f
C3024 avss.n56 dvss 0.18925f
C3025 avss.n57 dvss 0.115075f
C3026 avss.n58 dvss 0.218905f
C3027 avss.n59 dvss 0.151591f
C3028 avss.t313 dvss 1.38665f
C3029 avss.n60 dvss 0.636477f
C3030 avss.t19 dvss 0.315403f
C3031 avss.n61 dvss 0.201968f
C3032 avss.n62 dvss 0.228311f
C3033 avss.n63 dvss 0.855983f
C3034 avss.n64 dvss 0.133268f
C3035 avss.n65 dvss 0.855983f
C3036 avss.t109 dvss 7.42679f
C3037 avss.t300 dvss 0.273201f
C3038 avss.n66 dvss 1.75444f
C3039 avss.n67 dvss 55.1421f
C3040 avss.t312 dvss 9.758281f
C3041 avss.t224 dvss 11.6729f
C3042 avss.t139 dvss 11.6729f
C3043 avss.t220 dvss 11.6729f
C3044 avss.t101 dvss 11.5648f
C3045 avss.t177 dvss 11.6729f
C3046 avss.t221 dvss 11.6729f
C3047 avss.t194 dvss 11.6729f
C3048 avss.t222 dvss 11.6729f
C3049 avss.t200 dvss 11.6729f
C3050 avss.t191 dvss 11.6729f
C3051 avss.t193 dvss 11.6729f
C3052 avss.t116 dvss 11.6729f
C3053 avss.t253 dvss 11.6729f
C3054 avss.t255 dvss 5.94452f
C3055 avss.n68 dvss 68.3961f
C3056 avss.n69 dvss 40.7368f
C3057 avss.n117 dvss 0.812966f
C3058 avss.n128 dvss 0.337719f
C3059 avss.n129 dvss 0.332322f
C3060 avss.n140 dvss 0.337719f
C3061 avss.n141 dvss 0.332322f
C3062 avss.n152 dvss 0.337719f
C3063 avss.n153 dvss 0.332322f
C3064 avss.n164 dvss 0.337719f
C3065 avss.n165 dvss 0.332322f
C3066 avss.n176 dvss 0.337719f
C3067 avss.n177 dvss 0.332322f
C3068 avss.n188 dvss 0.337719f
C3069 avss.n189 dvss 0.332322f
C3070 avss.n200 dvss 0.337719f
C3071 avss.n201 dvss 0.332322f
C3072 avss.n212 dvss 0.337719f
C3073 avss.n213 dvss 0.332322f
C3074 avss.n224 dvss 0.337719f
C3075 avss.n225 dvss 0.332322f
C3076 avss.n236 dvss 0.337719f
C3077 avss.n237 dvss 0.332322f
C3078 avss.n248 dvss 0.337719f
C3079 avss.n249 dvss 0.332322f
C3080 avss.n260 dvss 0.337719f
C3081 avss.n261 dvss 0.332322f
C3082 avss.n272 dvss 0.337719f
C3083 avss.n273 dvss 0.332322f
C3084 avss.n284 dvss 0.337719f
C3085 avss.n285 dvss 0.332322f
C3086 avss.n296 dvss 0.337719f
C3087 avss.n297 dvss 0.332322f
C3088 avss.n307 dvss 0.408227f
C3089 avss.n308 dvss 13.633599f
C3090 avss.n320 dvss 0.216936f
C3091 avss.n321 dvss 6.86884f
C3092 avss.t271 dvss 10.0839f
C3093 avss.t122 dvss 10.0839f
C3094 avss.t205 dvss 10.0839f
C3095 avss.t104 dvss 10.0839f
C3096 avss.t123 dvss 10.0839f
C3097 avss.t335 dvss 10.0839f
C3098 avss.t251 dvss 10.0839f
C3099 avss.t105 dvss 10.604099f
C3100 avss.n322 dvss 5.76655f
C3101 avss.t213 dvss 5.21883f
C3102 avss.t83 dvss 0.315385f
C3103 avss.t77 dvss 0.315403f
C3104 avss.n323 dvss 0.195687f
C3105 avss.n324 dvss 0.188784f
C3106 avss.t73 dvss 0.315403f
C3107 avss.n325 dvss 0.195739f
C3108 avss.t79 dvss 0.315403f
C3109 avss.n326 dvss 0.193483f
C3110 avss.t75 dvss 0.315403f
C3111 avss.n327 dvss 0.193618f
C3112 avss.t51 dvss 0.315403f
C3113 avss.n328 dvss 0.19386f
C3114 avss.t29 dvss 0.315403f
C3115 avss.n329 dvss 0.157297f
C3116 avss.t7 dvss 0.315403f
C3117 avss.t21 dvss 0.315385f
C3118 avss.t31 dvss 0.315403f
C3119 avss.t11 dvss 0.315403f
C3120 avss.t64 dvss 0.315403f
C3121 avss.t27 dvss 0.315403f
C3122 avss.t55 dvss 0.315403f
C3123 avss.n330 dvss 0.202776f
C3124 avss.n331 dvss 0.193483f
C3125 avss.n332 dvss 0.193483f
C3126 avss.n333 dvss 0.193483f
C3127 avss.n334 dvss 0.195739f
C3128 avss.n335 dvss 0.188755f
C3129 avss.n336 dvss 0.192752f
C3130 avss.n338 dvss 0.255041f
C3131 avss.n339 dvss 0.289435f
C3132 avss.n340 dvss 0.863437f
C3133 avss.n341 dvss 5.83644f
C3134 avss.t258 dvss 3.44319f
C3135 avss.t279 dvss 5.52763f
C3136 avss.t280 dvss 3.05718f
C3137 avss.t178 dvss 2.74838f
C3138 avss.t56 dvss 5.18795f
C3139 avss.t187 dvss 3.39687f
C3140 avss.t130 dvss 2.74838f
C3141 avss.t188 dvss 4.84826f
C3142 avss.t28 dvss 3.73656f
C3143 avss.t156 dvss 2.74838f
C3144 avss.t135 dvss 2.91822f
C3145 avss.n342 dvss 2.74837f
C3146 avss.t136 dvss 2.91822f
C3147 avss.t257 dvss 2.74838f
C3148 avss.t65 dvss 4.16889f
C3149 avss.t334 dvss 4.41593f
C3150 avss.t128 dvss 2.74838f
C3151 avss.t331 dvss 3.8292f
C3152 avss.t12 dvss 4.75562f
C3153 avss.t103 dvss 2.74838f
C3154 avss.t327 dvss 3.48951f
C3155 avss.t328 dvss 5.09531f
C3156 avss.t336 dvss 2.74838f
C3157 avss.t32 dvss 3.14983f
C3158 avss.t155 dvss 5.43499f
C3159 avss.t208 dvss 2.74838f
C3160 avss.t152 dvss 2.81014f
C3161 avss.t22 dvss 5.49675f
C3162 avss.t182 dvss 3.0263f
C3163 avss.t192 dvss 2.74838f
C3164 avss.t183 dvss 5.21883f
C3165 avss.t8 dvss 3.36599f
C3166 avss.t102 dvss 2.74838f
C3167 avss.t365 dvss 4.87914f
C3168 avss.t362 dvss 3.70568f
C3169 avss.t119 dvss 2.74838f
C3170 avss.t30 dvss 4.53945f
C3171 avss.t289 dvss 4.04536f
C3172 avss.t250 dvss 2.74838f
C3173 avss.t288 dvss 4.19977f
C3174 avss.t52 dvss 4.38505f
C3175 avss.t129 dvss 2.74838f
C3176 avss.t325 dvss 3.86008f
C3177 avss.t322 dvss 4.72474f
C3178 avss.t272 dvss 2.74838f
C3179 avss.t76 dvss 3.52039f
C3180 avss.t162 dvss 5.06443f
C3181 avss.t176 dvss 2.74838f
C3182 avss.t161 dvss 3.18071f
C3183 avss.t80 dvss 5.40411f
C3184 avss.t0 dvss 2.74838f
C3185 avss.t131 dvss 2.84102f
C3186 avss.t134 dvss 5.49675f
C3187 avss.t74 dvss 2.99542f
C3188 avss.t310 dvss 2.74838f
C3189 avss.t219 dvss 5.24971f
C3190 avss.t216 dvss 3.33511f
C3191 avss.t157 dvss 2.74838f
C3192 avss.t84 dvss 4.91002f
C3193 avss.t112 dvss 3.6748f
C3194 avss.t249 dvss 2.74838f
C3195 avss.t113 dvss 4.57033f
C3196 avss.t78 dvss 4.01448f
C3197 avss.t214 dvss 2.74838f
C3198 avss.t273 dvss 4.23065f
C3199 avss.t274 dvss 4.35417f
C3200 avss.t215 dvss 2.74838f
C3201 avss.t20 dvss 3.89096f
C3202 avss.t306 dvss 4.69386f
C3203 avss.t341 dvss 2.74838f
C3204 avss.t305 dvss 4.24609f
C3205 avss.n343 dvss 5.03354f
C3206 avss.n344 dvss 0.863437f
C3207 avss.n346 dvss 0.260912f
C3208 avss.n348 dvss 1.10559f
C3209 avss.n349 dvss 3.13621f
C3210 avss.n350 dvss 0.718493f
C3211 avss.n351 dvss 1.43689f
C3212 avss.n352 dvss 1.28111f
C3213 avss.n353 dvss 1.09678f
C3214 avss.n354 dvss 0.61808f
C3215 avss.n355 dvss 3.90113f
C3216 avss.n356 dvss 0.850823f
C3217 avss.n357 dvss 0.411825f
C3218 avss.n358 dvss 0.979834f
C3219 avss.n359 dvss 0.802079f
C3220 avss.n360 dvss 0.79696f
C3221 avss.n361 dvss 0.79696f
C3222 avss.t16 dvss 0.151525p
C3223 avss.t108 dvss 16.6092f
C3224 avss.n362 dvss 3.34945f
C3225 avss.n363 dvss 30.546f
C3226 avss.t302 dvss 1.08873f
C3227 avss.n364 dvss 0.210762f
C3228 avss.n365 dvss 0.210762f
C3229 avss.t174 dvss 5.66035f
C3230 avss.t10 dvss 5.14638f
C3231 avss.n368 dvss 1.92787f
C3232 avss.n369 dvss 11.8829f
C3233 avss.n370 dvss 37.8865f
C3234 avss.n371 dvss 0.962219f
C3235 avss.n372 dvss 0.962219f
C3236 avss.n373 dvss 0.581746f
C3237 avss.n374 dvss 0.635632f
C3238 avss.n375 dvss 0.631795f
C3239 avss.n376 dvss 1.12119f
C3240 avss.t170 dvss 1.15678f
C3241 avss.n377 dvss 0.978815f
C3242 avss.t237 dvss 3.67895f
C3243 avss.t293 dvss 0.807024f
C3244 avss.n378 dvss 3.37863f
C3245 avss.t243 dvss 0.237245f
C3246 avss.t245 dvss 0.383655f
C3247 avss.t233 dvss 0.383655f
C3248 avss.t241 dvss 0.669852f
C3249 avss.n379 dvss 0.522874f
C3250 avss.n380 dvss 0.22497f
C3251 avss.n381 dvss 0.106394f
C3252 avss.n382 dvss 0.111001f
C3253 avss.n384 dvss 0.206591f
C3254 avss.n388 dvss 0.207128f
C3255 avss.n390 dvss 0.113335f
C3256 avss.n392 dvss 0.202403f
C3257 avss.n394 dvss 0.137583f
C3258 avss.n396 dvss 0.101505f
C3259 avss.n398 dvss 2.19514f
C3260 avss.n400 dvss 0.267313f
C3261 avss.n401 dvss 0.477684f
C3262 avss.t44 dvss 1.1347f
C3263 avss.t42 dvss 0.714783f
C3264 avss.n432 dvss 0.325671f
C3265 avss.n433 dvss 0.574646f
C3266 avss.n434 dvss 0.132287f
C3267 avss.n435 dvss 0.575305f
C3268 avss.n436 dvss 0.132188f
C3269 avss.n437 dvss 0.575305f
C3270 avss.n438 dvss 0.575305f
C3271 avss.n439 dvss 2.09896f
C3272 avss.n440 dvss 0.13249f
C3273 avss.n441 dvss 0.264395f
C3274 avss.n442 dvss 0.57554f
C3275 avss.n443 dvss 2.1139f
C3276 avss.n444 dvss 2.09896f
C3277 avss.n445 dvss 2.1139f
C3278 avss.n446 dvss 0.57554f
C3279 avss.n447 dvss 0.263987f
C3280 avss.n448 dvss 0.132187f
C3281 avss.n449 dvss 0.53745f
C3282 avss.n450 dvss 0.370954f
C3283 avss.n455 dvss 0.177133f
C3284 avss.n457 dvss 0.230764f
C3285 avss.t43 dvss 1.18286f
C3286 avss.n463 dvss 0.737479f
C3287 avss.n469 dvss 0.174096f
C3288 avss.n473 dvss 1.57797f
C3289 avss.n477 dvss 0.177133f
C3290 avss.n480 dvss 0.240951f
C3291 avss.n482 dvss 0.240951f
C3292 avss.n488 dvss 0.177133f
C3293 avss.n489 dvss 0.793494f
C3294 avss.n496 dvss 0.236822f
C3295 avss.n497 dvss 0.236822f
C3296 avss.n498 dvss 0.174096f
C3297 avss.n505 dvss 0.761839f
C3298 avss.n506 dvss 0.226632f
C3299 avss.n507 dvss 1.46802f
C3300 avss.n513 dvss 0.226632f
C3301 avss.n514 dvss 1.44122f
C3302 avss.n522 dvss 0.169643f
C3303 avss.n523 dvss 0.169643f
C3304 avss.n524 dvss 0.230764f
C3305 avss.n530 dvss 1.52357f
C3306 avss.n531 dvss 0.784423f
C3307 avss.n532 dvss 0.177133f
C3308 avss.n536 dvss 0.121899f
C3309 avss.n537 dvss 3.79452f
C3310 avss.n538 dvss 14.446599f
C3311 avss.t380 dvss 1.75819f
C3312 avss.n539 dvss 1.73465f
C3313 avss.t60 dvss 1.1347f
C3314 avss.n540 dvss 0.56215f
C3315 avss.n542 dvss 0.477684f
C3316 avss.n544 dvss 0.137583f
C3317 avss.n546 dvss 0.127047f
C3318 avss.n547 dvss 0.476407f
C3319 avss.n548 dvss 1.1811f
C3320 avss.n550 dvss 0.102779f
C3321 avss.n551 dvss 0.476407f
C3322 avss.n552 dvss 0.581746f
C3323 avss.n553 dvss 0.953696f
C3324 avss.n556 dvss 0.126186f
C3325 avss.n557 dvss 0.216416f
C3326 avss.n558 dvss 0.216416f
C3327 avss.t295 dvss 2.16927f
C3328 avss.n560 dvss 0.124229f
C3329 avss.n561 dvss 0.210762f
C3330 avss.n562 dvss 2.89614f
C3331 avss.t360 dvss 1.2419f
C3332 avss.t311 dvss 11.819401f
C3333 avss.n563 dvss 0.797033f
C3334 avss.t264 dvss 11.3332f
C3335 avss.t195 dvss 14.1384f
C3336 avss.t287 dvss 14.1384f
C3337 avss.t309 dvss 14.1384f
C3338 avss.t106 dvss 10.6038f
C3339 avss.t263 dvss 14.1384f
C3340 avss.t118 dvss 14.1384f
C3341 avss.t207 dvss 14.1384f
C3342 avss.t223 dvss 14.1384f
C3343 avss.t184 dvss 14.1384f
C3344 avss.t303 dvss 14.1384f
C3345 avss.t107 dvss 14.1384f
C3346 avss.t140 dvss 14.1384f
C3347 avss.t117 dvss 10.6038f
C3348 avss.n564 dvss 7.06922f
C3349 avss.n565 dvss 0.797033f
C3350 avss.n566 dvss 0.400895f
C3351 avss.n567 dvss 0.676991f
C3352 avss.t259 dvss 9.87447f
C3353 avss.t150 dvss 14.1384f
C3354 avss.t100 dvss 14.1384f
C3355 avss.t202 dvss 14.1384f
C3356 avss.t321 dvss 13.8082f
C3357 avss.n568 dvss 35.874897f
C3358 avss.n569 dvss 0.794576f
C3359 avss.n571 dvss 0.206591f
C3360 avss.n575 dvss 0.207128f
C3361 avss.n577 dvss 0.113335f
C3362 avss.n579 dvss 0.115437f
C3363 avss.n580 dvss 0.111001f
C3364 avss.n581 dvss 0.131177f
C3365 avss.n582 dvss 0.522874f
C3366 avss.n583 dvss 1.01798f
C3367 avss.t356 dvss 0.669852f
C3368 avss.t346 dvss 0.383655f
C3369 avss.t350 dvss 0.383655f
C3370 avss.t352 dvss 0.383655f
C3371 avss.t344 dvss 0.287738f
C3372 avss.n584 dvss 0.195137f
C3373 avss.n585 dvss 0.105949f
C3374 avss.n587 dvss 0.21913f
C3375 avss.n588 dvss 0.112073f
C3376 avss.t40 dvss 7.17465f
C3377 avss.n589 dvss 0.962219f
C3378 avss.n590 dvss 0.301526f
C3379 avss.n591 dvss 0.267313f
C3380 avss.n592 dvss 0.127047f
C3381 avss.t39 dvss 1.1347f
C3382 avss.n593 dvss 0.267313f
C3383 avss.t46 dvss 1.1347f
C3384 avss.n596 dvss 0.56215f
C3385 avss.t387 dvss 1.75819f
C3386 avss.n598 dvss 0.807458f
C3387 avss.t366 dvss 1.75819f
C3388 avss.n599 dvss 0.807458f
C3389 avss.t377 dvss 1.75819f
C3390 avss.n600 dvss 0.807458f
C3391 avss.t397 dvss 1.75819f
C3392 avss.n601 dvss 0.807458f
C3393 avss.t375 dvss 1.75819f
C3394 avss.n602 dvss 0.807458f
C3395 avss.t382 dvss 1.75819f
C3396 avss.n603 dvss 0.807458f
C3397 avss.t393 dvss 1.75819f
C3398 avss.n604 dvss 0.892742f
C3399 avss.n605 dvss 0.220039f
C3400 avss.n607 dvss 0.56215f
C3401 avss.n609 dvss 0.137583f
C3402 avss.n610 dvss 0.477684f
C3403 avss.n612 dvss 0.138274f
C3404 avss.n613 dvss 0.635632f
C3405 avss.n614 dvss 0.547309f
C3406 avss.t229 dvss 9.07712f
C3407 avss.t227 dvss 6.80784f
C3408 avss.t61 dvss 7.17465f
C3409 avss.t231 dvss 9.07712f
C3410 avss.t225 dvss 6.80784f
C3411 avss.n615 dvss 4.53856f
C3412 avss.n616 dvss 0.953696f
C3413 avss.n617 dvss 0.962219f
C3414 avss.n618 dvss 3.02007f
C3415 avss.n619 dvss 0.248186f
C3416 avss.t358 dvss 0.291727f
C3417 avss.t342 dvss 0.383655f
C3418 avss.t354 dvss 0.383655f
C3419 avss.t348 dvss 0.287738f
C3420 avss.n621 dvss 0.21913f
C3421 avss.n623 dvss 0.105949f
C3422 avss.n624 dvss 0.283477f
C3423 avss.n625 dvss 0.581378f
C3424 avss.n626 dvss 0.398522f
C3425 avss.n627 dvss 0.936463f
C3426 avss.n628 dvss 1.09871f
C3427 avss.n629 dvss 1.07854f
C3428 avss.n630 dvss 0.797033f
C3429 avss.n631 dvss 0.79696f
C3430 avss.n632 dvss 0.79696f
C3431 avss.n633 dvss 11.6698f
C3432 avss.t297 dvss 2.06733f
C3433 avss.n634 dvss 33.297302f
C3434 avss.n635 dvss 29.9021f
C3435 avss.t14 dvss 23.9296f
C3436 avss.n636 dvss 0.664573f
C3437 avss.n637 dvss 0.664573f
C3438 avss.n638 dvss 0.206801f
C3439 avss.n639 dvss 0.206801f
C3440 avss.n640 dvss 0.693973f
C3441 avss.n641 dvss 0.357435f
C3442 avss.t69 dvss 0.156831f
C3443 avss.t68 dvss 1.84402f
C3444 avss.n642 dvss 1.633f
C3445 avss.n643 dvss 0.716895f
C3446 avss.t13 dvss 2.3615f
C3447 avss.n644 dvss 1.8839f
C3448 avss.t36 dvss 0.156831f
C3449 avss.t35 dvss 1.84402f
C3450 avss.n645 dvss 1.633f
C3451 avss.n646 dvss 0.718878f
C3452 avss.n647 dvss 0.502253f
C3453 avss.n648 dvss 0.2001f
C3454 avss.n649 dvss 0.2001f
C3455 avss.t114 dvss 4.97584f
C3456 avss.t282 dvss 6.10827f
C3457 avss.t281 dvss 6.10827f
C3458 avss.n650 dvss 0.406171f
C3459 avss.t115 dvss 51.6545f
C3460 avss.n652 dvss 0.400092f
C3461 avss.n653 dvss 0.411825f
C3462 avss.n654 dvss 0.811972f
C3463 avss.n655 dvss 0.716607f
C3464 avss.t209 dvss 0.237267f
C3465 avss.n656 dvss 1.09388f
C3466 avss.n657 dvss 0.724867f
C3467 avss.n658 dvss 0.714341f
C3468 avss.n659 dvss 0.598349f
C3469 avss.n660 dvss 0.797033f
C3470 avss.n661 dvss 22.5139f
C3471 avss.n662 dvss 17.058f
C3472 avss.n663 dvss 0.658058f
C3473 avss.n664 dvss 0.386557f
C3474 avss.n665 dvss 0.673184f
C3475 avss.n666 dvss 0.693973f
C3476 avss.n667 dvss 0.637517f
C3477 avss.n668 dvss 0.373176f
C3478 avss.n669 dvss 0.658058f
C3479 avss.n670 dvss 24.155699f
C3480 avss.n671 dvss 31.2904f
C3481 avss.n672 dvss 16.009201f
C3482 avss.t267 dvss 0.809095f
C3483 avss.n673 dvss 1.39406f
C3484 avss.t269 dvss 2.19475f
C3485 avss.t265 dvss 1.23275f
C3486 avss.n674 dvss 1.13401f
C3487 avss.n675 dvss 0.210762f
C3488 avss.n678 dvss 0.301526f
C3489 avss.n679 dvss 0.547309f
C3490 avss.n680 dvss 0.631795f
C3491 avss.n682 dvss 2.19514f
C3492 avss.n683 dvss 0.212919f
C3493 avss.n684 dvss 0.102174f
C3494 avss.n685 dvss 0.11336f
C3495 avss.n686 dvss 0.315931f
C3496 avss.n687 dvss 1.26368f
C3497 avss.t70 dvss 1.1347f
C3498 avss.n688 dvss 0.56215f
C3499 avss.n691 dvss 0.267313f
C3500 avss.n692 dvss 0.267313f
C3501 avss.n693 dvss 0.222831f
C3502 avss.t383 dvss 1.74585f
C3503 avss.n694 dvss 0.884212f
C3504 avss.t372 dvss 1.74585f
C3505 avss.n695 dvss 0.792955f
C3506 avss.t367 dvss 1.74585f
C3507 avss.n696 dvss 0.792955f
C3508 avss.t389 dvss 1.74585f
C3509 avss.n697 dvss 0.792955f
C3510 avss.t368 dvss 1.74585f
C3511 avss.n698 dvss 0.792955f
C3512 avss.t390 dvss 1.74585f
C3513 avss.n699 dvss 0.792955f
C3514 avss.t373 dvss 1.74585f
C3515 avss.n700 dvss 0.792955f
C3516 avss.t371 dvss 1.74585f
C3517 avss.n701 dvss 0.846411f
C3518 avss.n702 dvss 4.00717f
C3519 avss.n703 dvss 11.1399f
C3520 avss.n704 dvss 13.7076f
C3521 avss.n705 dvss 10.085401f
C3522 avss.t23 dvss 1.1347f
C3523 avss.n706 dvss 0.56215f
C3524 avss.n708 dvss 0.477684f
C3525 avss.n710 dvss 0.137583f
C3526 avss.n712 dvss 0.127047f
C3527 avss.n713 dvss 0.476407f
C3528 avss.n714 dvss 0.212919f
C3529 avss.n715 dvss 0.102174f
C3530 avss.n716 dvss 0.11336f
C3531 avss.n717 dvss 0.383744f
C3532 avss.n718 dvss 1.26368f
C3533 avss.t85 dvss 1.1347f
C3534 avss.n719 dvss 0.56215f
C3535 avss.n722 dvss 0.267313f
C3536 avss.n723 dvss 0.267313f
C3537 avss.n724 dvss 0.222831f
C3538 avss.t388 dvss 1.74585f
C3539 avss.n725 dvss 0.884212f
C3540 avss.t391 dvss 1.74585f
C3541 avss.n726 dvss 0.792955f
C3542 avss.t395 dvss 1.74585f
C3543 avss.n727 dvss 0.792955f
C3544 avss.t378 dvss 1.74585f
C3545 avss.n728 dvss 0.792955f
C3546 avss.t394 dvss 1.74585f
C3547 avss.n729 dvss 0.792955f
C3548 avss.t370 dvss 1.74585f
C3549 avss.n730 dvss 0.792955f
C3550 avss.t385 dvss 1.74585f
C3551 avss.n731 dvss 0.792955f
C3552 avss.t392 dvss 1.74585f
C3553 avss.n732 dvss 0.846411f
C3554 avss.n733 dvss 6.9307f
C3555 avss.t381 dvss 1.75819f
C3556 avss.n734 dvss 1.73465f
C3557 avss.t374 dvss 1.75819f
C3558 avss.n735 dvss 0.807458f
C3559 avss.t396 dvss 1.75819f
C3560 avss.n736 dvss 0.807458f
C3561 avss.t384 dvss 1.75819f
C3562 avss.n737 dvss 0.807458f
C3563 avss.t369 dvss 1.75819f
C3564 avss.n738 dvss 0.807458f
C3565 avss.t386 dvss 1.75819f
C3566 avss.n739 dvss 0.807458f
C3567 avss.t379 dvss 1.75819f
C3568 avss.n740 dvss 0.807458f
C3569 avss.t376 dvss 1.75819f
C3570 avss.n741 dvss 0.892742f
C3571 avss.n742 dvss 0.220039f
C3572 avss.n744 dvss 0.56215f
C3573 avss.n746 dvss 0.137583f
C3574 avss.t1 dvss 1.1347f
C3575 avss.n747 dvss 0.56215f
C3576 avss.n749 dvss 0.127047f
C3577 avss.n750 dvss 0.476407f
C3578 avss.n751 dvss 0.267313f
C3579 avss.n753 dvss 1.1811f
C3580 avss.n754 dvss 0.195137f
C3581 avss.n755 dvss 0.105949f
C3582 avss.n756 dvss 0.21913f
C3583 avss.n758 dvss 0.131177f
C3584 avss.n760 dvss 0.21913f
C3585 avss.t24 dvss 2.59831f
C3586 avss.n762 dvss 0.615877f
C3587 avss.t172 dvss 3.79677f
C3588 avss.n763 dvss 3.1678f
C3589 avss.t235 dvss 2.74604f
C3590 avss.t2 dvss 3.1678f
C3591 avss.t239 dvss 4.30612f
C3592 avss.t247 dvss 4.35522f
C3593 avss.n765 dvss 1.5839f
C3594 avss.n766 dvss 0.953696f
C3595 avss.n767 dvss 0.547309f
C3596 avss.n769 dvss 0.301526f
C3597 avss.n771 dvss 0.301526f
C3598 avss.n772 dvss 0.547309f
C3599 avss.n773 dvss 0.953696f
C3600 avss.n774 dvss 3.96865f
C3601 avss.n775 dvss 0.216416f
C3602 avss.n777 dvss 0.124229f
C3603 avss.n778 dvss 0.126186f
C3604 avss.n779 dvss 0.216416f
C3605 avss.n780 dvss 4.41173f
C3606 avss.n781 dvss 35.307602f
C3607 avss.n782 dvss 39.4683f
C3608 avss.n783 dvss 0.797033f
C3609 avss.n784 dvss 0.592037f
C3610 avss.n785 dvss 0.687297f
C3611 avss.n786 dvss 0.786545f
C3612 avss.n787 dvss 0.743352f
C3613 avss.n788 dvss 7.84116f
C3614 avss.n789 dvss 4.872221f
C3615 avss.n790 dvss 0.134145f
C3616 avss.n791 dvss 1.53113f
C3617 avss.n792 dvss 1.54882f
C3618 avss.n793 dvss 2.89223f
C3619 avss.n794 dvss 2.88571f
C3620 avss.n795 dvss 1.75259f
C3621 avss.n796 dvss 1.75444f
C3622 avss.n797 dvss 1.75444f
C3623 avss.n798 dvss 1.68985f
C3624 avss.t143 dvss -1.14557f
C3625 avss.t82 dvss 5.19758f
C3626 avss.t185 dvss 4.55749f
C3627 avss.t320 dvss 6.78502f
C3628 avss.t54 dvss 7.45073f
C3629 avss.t99 dvss 4.55749f
C3630 avss.t319 dvss 6.22174f
C3631 avss.t292 dvss 4.68551f
C3632 avss.n799 dvss 0.654931f
C3633 avss.n800 dvss 1.10882f
C3634 avss.n801 dvss 3.45652f
C3635 avss.n802 dvss 1.10882f
C3636 avss.n803 dvss 0.653173f
C3637 avss.n804 dvss 0.756922f
C3638 avss.n805 dvss 0.165885f
C3639 avss.n806 dvss 1.27521f
C3640 avss.n807 dvss 1.27521f
C3641 avss.t66 dvss 4.16156f
C3642 avss.n808 dvss 0.165885f
C3643 avss.t67 dvss 0.204737f
C3644 avss.n809 dvss 1.57106f
C3645 avss.n810 dvss 0.466083f
C3646 avss.n811 dvss 0.201653f
C3647 avss.n812 dvss 0.510971f
C3648 avss.n813 dvss 0.466083f
C3649 avss.t33 dvss 4.16156f
C3650 avss.n814 dvss 1.57106f
C3651 avss.t34 dvss 0.204737f
C3652 avss.n815 dvss 0.165885f
C3653 avss.n816 dvss 1.27521f
C3654 avss.n817 dvss 0.165885f
C3655 avss.n818 dvss 1.27521f
C3656 avss.t57 dvss 4.16156f
C3657 avss.t59 dvss 0.16157f
C3658 avss.n819 dvss 1.57106f
C3659 avss.n820 dvss 0.407738f
C3660 avss.n821 dvss 0.275557f
C3661 avss.n822 dvss 0.510532f
C3662 avss.n823 dvss 0.201214f
C3663 avss.n824 dvss 0.275557f
C3664 avss.n825 dvss 1.04504f
C3665 avss.n826 dvss 1.04504f
C3666 avss.n827 dvss 0.275557f
C3667 avss.t93 dvss 4.16156f
C3668 avss.t95 dvss 0.16157f
C3669 avss.n828 dvss 1.57106f
C3670 avss.n829 dvss 0.407738f
C3671 avss.n830 dvss 0.165885f
C3672 avss.n831 dvss 1.27521f
C3673 avss.n832 dvss 1.27521f
C3674 avss.t4 dvss 4.16156f
C3675 avss.n833 dvss 0.165885f
C3676 avss.t6 dvss 0.204737f
C3677 avss.n834 dvss 1.57106f
C3678 avss.n835 dvss 0.466083f
C3679 avss.n836 dvss 0.153927f
C3680 avss.n837 dvss 0.226735f
C3681 avss.n838 dvss 0.466083f
C3682 avss.t96 dvss 4.16156f
C3683 avss.n839 dvss 1.57106f
C3684 avss.t97 dvss 0.204737f
C3685 avss.n840 dvss 0.165885f
C3686 avss.n841 dvss 1.27521f
C3687 avss.n842 dvss 0.165885f
C3688 avss.n843 dvss 1.27521f
C3689 avss.t90 dvss 4.16156f
C3690 avss.t92 dvss 0.16157f
C3691 avss.n844 dvss 1.57106f
C3692 avss.n845 dvss 0.407738f
C3693 avss.n846 dvss 0.275557f
C3694 avss.n847 dvss 0.226296f
C3695 avss.n848 dvss 0.458673f
C3696 avss.n849 dvss 0.275557f
C3697 avss.n850 dvss 1.06482f
C3698 avss.n851 dvss 1.1042f
C3699 avss.n852 dvss 0.873523f
C3700 avss.n853 dvss 0.152472f
C3701 avss.n854 dvss 0.20668f
C3702 avss.n855 dvss 0.152472f
C3703 avss.n856 dvss 0.131025f
C3704 avss.n857 dvss 0.406171f
C3705 avss.n858 dvss 6.52899f
C3706 avss.n859 dvss 7.42512f
C3707 avss.n860 dvss 0.302087f
C3708 avss.n861 dvss 0.100638f
C3709 avss.n862 dvss 0.122092f
C3710 avss.n863 dvss 0.111751f
C3711 avss.t197 dvss 0.216631f
C3712 avss.n864 dvss 0.425304f
C3713 avss.n865 dvss 0.158735f
C3714 avss.n866 dvss 0.569362f
C3715 avss.t318 dvss 0.216631f
C3716 avss.n867 dvss 0.425524f
C3717 avss.n868 dvss 0.157574f
C3718 avss.n869 dvss 0.122092f
C3719 avss.n870 dvss 0.100638f
C3720 avss.n871 dvss 0.302087f
C3721 avss.n872 dvss 2.27874f
C3722 avss.t5 dvss 6.17053f
C3723 avss.n873 dvss 7.39952f
C3724 avss.n874 dvss 0.209014f
C3725 avss.n875 dvss 0.115267f
C3726 avss.n876 dvss 0.304253f
C3727 avss.n877 dvss 0.115773f
C3728 avss.n878 dvss 0.209014f
C3729 avss.n879 dvss 9.67826f
C3730 avss.t314 dvss 13.314f
C3731 avss.t212 dvss 10.9072f
C3732 avss.n880 dvss 20.613598f
C3733 avss.t167 dvss 17.8407f
C3734 avss.t210 dvss 15.683701f
C3735 avss.t206 dvss 15.826401f
C3736 avss.t211 dvss 15.826401f
C3737 avss.t98 dvss 15.826401f
C3738 avss.t203 dvss 15.826401f
C3739 avss.t256 dvss 12.7072f
C3740 avss.n881 dvss 17.7825f
C3741 avss.n882 dvss 12.4021f
C3742 avss.t120 dvss 2.8022f
C3743 avss.n888 dvss 0.159932f
C3744 avss.n889 dvss 0.336259f
C3745 avss.n890 dvss 0.575862f
C3746 avss.n891 dvss 0.426899f
.ends


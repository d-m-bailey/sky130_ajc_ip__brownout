magic
tech sky130A
magscale 1 2
timestamp 1712590844
<< nwell >>
rect -5203 -909 5203 909
<< mvpmos >>
rect -4945 483 -3345 683
rect -3287 483 -1687 683
rect -1629 483 -29 683
rect 29 483 1629 683
rect 1687 483 3287 683
rect 3345 483 4945 683
rect -4945 118 -3345 318
rect -3287 118 -1687 318
rect -1629 118 -29 318
rect 29 118 1629 318
rect 1687 118 3287 318
rect 3345 118 4945 318
rect -4945 -247 -3345 -47
rect -3287 -247 -1687 -47
rect -1629 -247 -29 -47
rect 29 -247 1629 -47
rect 1687 -247 3287 -47
rect 3345 -247 4945 -47
rect -4945 -612 -3345 -412
rect -3287 -612 -1687 -412
rect -1629 -612 -29 -412
rect 29 -612 1629 -412
rect 1687 -612 3287 -412
rect 3345 -612 4945 -412
<< mvpdiff >>
rect -5003 671 -4945 683
rect -5003 495 -4991 671
rect -4957 495 -4945 671
rect -5003 483 -4945 495
rect -3345 671 -3287 683
rect -3345 495 -3333 671
rect -3299 495 -3287 671
rect -3345 483 -3287 495
rect -1687 671 -1629 683
rect -1687 495 -1675 671
rect -1641 495 -1629 671
rect -1687 483 -1629 495
rect -29 671 29 683
rect -29 495 -17 671
rect 17 495 29 671
rect -29 483 29 495
rect 1629 671 1687 683
rect 1629 495 1641 671
rect 1675 495 1687 671
rect 1629 483 1687 495
rect 3287 671 3345 683
rect 3287 495 3299 671
rect 3333 495 3345 671
rect 3287 483 3345 495
rect 4945 671 5003 683
rect 4945 495 4957 671
rect 4991 495 5003 671
rect 4945 483 5003 495
rect -5003 306 -4945 318
rect -5003 130 -4991 306
rect -4957 130 -4945 306
rect -5003 118 -4945 130
rect -3345 306 -3287 318
rect -3345 130 -3333 306
rect -3299 130 -3287 306
rect -3345 118 -3287 130
rect -1687 306 -1629 318
rect -1687 130 -1675 306
rect -1641 130 -1629 306
rect -1687 118 -1629 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 1629 306 1687 318
rect 1629 130 1641 306
rect 1675 130 1687 306
rect 1629 118 1687 130
rect 3287 306 3345 318
rect 3287 130 3299 306
rect 3333 130 3345 306
rect 3287 118 3345 130
rect 4945 306 5003 318
rect 4945 130 4957 306
rect 4991 130 5003 306
rect 4945 118 5003 130
rect -5003 -59 -4945 -47
rect -5003 -235 -4991 -59
rect -4957 -235 -4945 -59
rect -5003 -247 -4945 -235
rect -3345 -59 -3287 -47
rect -3345 -235 -3333 -59
rect -3299 -235 -3287 -59
rect -3345 -247 -3287 -235
rect -1687 -59 -1629 -47
rect -1687 -235 -1675 -59
rect -1641 -235 -1629 -59
rect -1687 -247 -1629 -235
rect -29 -59 29 -47
rect -29 -235 -17 -59
rect 17 -235 29 -59
rect -29 -247 29 -235
rect 1629 -59 1687 -47
rect 1629 -235 1641 -59
rect 1675 -235 1687 -59
rect 1629 -247 1687 -235
rect 3287 -59 3345 -47
rect 3287 -235 3299 -59
rect 3333 -235 3345 -59
rect 3287 -247 3345 -235
rect 4945 -59 5003 -47
rect 4945 -235 4957 -59
rect 4991 -235 5003 -59
rect 4945 -247 5003 -235
rect -5003 -424 -4945 -412
rect -5003 -600 -4991 -424
rect -4957 -600 -4945 -424
rect -5003 -612 -4945 -600
rect -3345 -424 -3287 -412
rect -3345 -600 -3333 -424
rect -3299 -600 -3287 -424
rect -3345 -612 -3287 -600
rect -1687 -424 -1629 -412
rect -1687 -600 -1675 -424
rect -1641 -600 -1629 -424
rect -1687 -612 -1629 -600
rect -29 -424 29 -412
rect -29 -600 -17 -424
rect 17 -600 29 -424
rect -29 -612 29 -600
rect 1629 -424 1687 -412
rect 1629 -600 1641 -424
rect 1675 -600 1687 -424
rect 1629 -612 1687 -600
rect 3287 -424 3345 -412
rect 3287 -600 3299 -424
rect 3333 -600 3345 -424
rect 3287 -612 3345 -600
rect 4945 -424 5003 -412
rect 4945 -600 4957 -424
rect 4991 -600 5003 -424
rect 4945 -612 5003 -600
<< mvpdiffc >>
rect -4991 495 -4957 671
rect -3333 495 -3299 671
rect -1675 495 -1641 671
rect -17 495 17 671
rect 1641 495 1675 671
rect 3299 495 3333 671
rect 4957 495 4991 671
rect -4991 130 -4957 306
rect -3333 130 -3299 306
rect -1675 130 -1641 306
rect -17 130 17 306
rect 1641 130 1675 306
rect 3299 130 3333 306
rect 4957 130 4991 306
rect -4991 -235 -4957 -59
rect -3333 -235 -3299 -59
rect -1675 -235 -1641 -59
rect -17 -235 17 -59
rect 1641 -235 1675 -59
rect 3299 -235 3333 -59
rect 4957 -235 4991 -59
rect -4991 -600 -4957 -424
rect -3333 -600 -3299 -424
rect -1675 -600 -1641 -424
rect -17 -600 17 -424
rect 1641 -600 1675 -424
rect 3299 -600 3333 -424
rect 4957 -600 4991 -424
<< mvnsubdiff >>
rect -5137 831 5137 843
rect -5137 797 -5029 831
rect 5029 797 5137 831
rect -5137 785 5137 797
rect -5137 735 -5079 785
rect -5137 -735 -5125 735
rect -5091 -735 -5079 735
rect 5079 735 5137 785
rect -5137 -785 -5079 -735
rect 5079 -735 5091 735
rect 5125 -735 5137 735
rect 5079 -785 5137 -735
rect -5137 -797 5137 -785
rect -5137 -831 -5029 -797
rect 5029 -831 5137 -797
rect -5137 -843 5137 -831
<< mvnsubdiffcont >>
rect -5029 797 5029 831
rect -5125 -735 -5091 735
rect 5091 -735 5125 735
rect -5029 -831 5029 -797
<< poly >>
rect -4945 683 -3345 709
rect -3287 683 -1687 709
rect -1629 683 -29 709
rect 29 683 1629 709
rect 1687 683 3287 709
rect 3345 683 4945 709
rect -4945 436 -3345 483
rect -4945 402 -4929 436
rect -3361 402 -3345 436
rect -4945 386 -3345 402
rect -3287 436 -1687 483
rect -3287 402 -3271 436
rect -1703 402 -1687 436
rect -3287 386 -1687 402
rect -1629 436 -29 483
rect -1629 402 -1613 436
rect -45 402 -29 436
rect -1629 386 -29 402
rect 29 436 1629 483
rect 29 402 45 436
rect 1613 402 1629 436
rect 29 386 1629 402
rect 1687 436 3287 483
rect 1687 402 1703 436
rect 3271 402 3287 436
rect 1687 386 3287 402
rect 3345 436 4945 483
rect 3345 402 3361 436
rect 4929 402 4945 436
rect 3345 386 4945 402
rect -4945 318 -3345 344
rect -3287 318 -1687 344
rect -1629 318 -29 344
rect 29 318 1629 344
rect 1687 318 3287 344
rect 3345 318 4945 344
rect -4945 71 -3345 118
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -4945 21 -3345 37
rect -3287 71 -1687 118
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -3287 21 -1687 37
rect -1629 71 -29 118
rect -1629 37 -1613 71
rect -45 37 -29 71
rect -1629 21 -29 37
rect 29 71 1629 118
rect 29 37 45 71
rect 1613 37 1629 71
rect 29 21 1629 37
rect 1687 71 3287 118
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 1687 21 3287 37
rect 3345 71 4945 118
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 3345 21 4945 37
rect -4945 -47 -3345 -21
rect -3287 -47 -1687 -21
rect -1629 -47 -29 -21
rect 29 -47 1629 -21
rect 1687 -47 3287 -21
rect 3345 -47 4945 -21
rect -4945 -294 -3345 -247
rect -4945 -328 -4929 -294
rect -3361 -328 -3345 -294
rect -4945 -344 -3345 -328
rect -3287 -294 -1687 -247
rect -3287 -328 -3271 -294
rect -1703 -328 -1687 -294
rect -3287 -344 -1687 -328
rect -1629 -294 -29 -247
rect -1629 -328 -1613 -294
rect -45 -328 -29 -294
rect -1629 -344 -29 -328
rect 29 -294 1629 -247
rect 29 -328 45 -294
rect 1613 -328 1629 -294
rect 29 -344 1629 -328
rect 1687 -294 3287 -247
rect 1687 -328 1703 -294
rect 3271 -328 3287 -294
rect 1687 -344 3287 -328
rect 3345 -294 4945 -247
rect 3345 -328 3361 -294
rect 4929 -328 4945 -294
rect 3345 -344 4945 -328
rect -4945 -412 -3345 -386
rect -3287 -412 -1687 -386
rect -1629 -412 -29 -386
rect 29 -412 1629 -386
rect 1687 -412 3287 -386
rect 3345 -412 4945 -386
rect -4945 -659 -3345 -612
rect -4945 -693 -4929 -659
rect -3361 -693 -3345 -659
rect -4945 -709 -3345 -693
rect -3287 -659 -1687 -612
rect -3287 -693 -3271 -659
rect -1703 -693 -1687 -659
rect -3287 -709 -1687 -693
rect -1629 -659 -29 -612
rect -1629 -693 -1613 -659
rect -45 -693 -29 -659
rect -1629 -709 -29 -693
rect 29 -659 1629 -612
rect 29 -693 45 -659
rect 1613 -693 1629 -659
rect 29 -709 1629 -693
rect 1687 -659 3287 -612
rect 1687 -693 1703 -659
rect 3271 -693 3287 -659
rect 1687 -709 3287 -693
rect 3345 -659 4945 -612
rect 3345 -693 3361 -659
rect 4929 -693 4945 -659
rect 3345 -709 4945 -693
<< polycont >>
rect -4929 402 -3361 436
rect -3271 402 -1703 436
rect -1613 402 -45 436
rect 45 402 1613 436
rect 1703 402 3271 436
rect 3361 402 4929 436
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect -4929 -328 -3361 -294
rect -3271 -328 -1703 -294
rect -1613 -328 -45 -294
rect 45 -328 1613 -294
rect 1703 -328 3271 -294
rect 3361 -328 4929 -294
rect -4929 -693 -3361 -659
rect -3271 -693 -1703 -659
rect -1613 -693 -45 -659
rect 45 -693 1613 -659
rect 1703 -693 3271 -659
rect 3361 -693 4929 -659
<< locali >>
rect -5125 797 -5029 831
rect 5029 797 5125 831
rect -5125 735 -5091 797
rect 5091 735 5125 797
rect -4991 671 -4957 687
rect -4991 479 -4957 495
rect -3333 671 -3299 687
rect -3333 479 -3299 495
rect -1675 671 -1641 687
rect -1675 479 -1641 495
rect -17 671 17 687
rect -17 479 17 495
rect 1641 671 1675 687
rect 1641 479 1675 495
rect 3299 671 3333 687
rect 3299 479 3333 495
rect 4957 671 4991 687
rect 4957 479 4991 495
rect -4945 402 -4929 436
rect -3361 402 -3345 436
rect -3287 402 -3271 436
rect -1703 402 -1687 436
rect -1629 402 -1613 436
rect -45 402 -29 436
rect 29 402 45 436
rect 1613 402 1629 436
rect 1687 402 1703 436
rect 3271 402 3287 436
rect 3345 402 3361 436
rect 4929 402 4945 436
rect -4991 306 -4957 322
rect -4991 114 -4957 130
rect -3333 306 -3299 322
rect -3333 114 -3299 130
rect -1675 306 -1641 322
rect -1675 114 -1641 130
rect -17 306 17 322
rect -17 114 17 130
rect 1641 306 1675 322
rect 1641 114 1675 130
rect 3299 306 3333 322
rect 3299 114 3333 130
rect 4957 306 4991 322
rect 4957 114 4991 130
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -1629 37 -1613 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1613 37 1629 71
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 3345 37 3361 71
rect 4929 37 4945 71
rect -4991 -59 -4957 -43
rect -4991 -251 -4957 -235
rect -3333 -59 -3299 -43
rect -3333 -251 -3299 -235
rect -1675 -59 -1641 -43
rect -1675 -251 -1641 -235
rect -17 -59 17 -43
rect -17 -251 17 -235
rect 1641 -59 1675 -43
rect 1641 -251 1675 -235
rect 3299 -59 3333 -43
rect 3299 -251 3333 -235
rect 4957 -59 4991 -43
rect 4957 -251 4991 -235
rect -4945 -328 -4929 -294
rect -3361 -328 -3345 -294
rect -3287 -328 -3271 -294
rect -1703 -328 -1687 -294
rect -1629 -328 -1613 -294
rect -45 -328 -29 -294
rect 29 -328 45 -294
rect 1613 -328 1629 -294
rect 1687 -328 1703 -294
rect 3271 -328 3287 -294
rect 3345 -328 3361 -294
rect 4929 -328 4945 -294
rect -4991 -424 -4957 -408
rect -4991 -616 -4957 -600
rect -3333 -424 -3299 -408
rect -3333 -616 -3299 -600
rect -1675 -424 -1641 -408
rect -1675 -616 -1641 -600
rect -17 -424 17 -408
rect -17 -616 17 -600
rect 1641 -424 1675 -408
rect 1641 -616 1675 -600
rect 3299 -424 3333 -408
rect 3299 -616 3333 -600
rect 4957 -424 4991 -408
rect 4957 -616 4991 -600
rect -4945 -693 -4929 -659
rect -3361 -693 -3345 -659
rect -3287 -693 -3271 -659
rect -1703 -693 -1687 -659
rect -1629 -693 -1613 -659
rect -45 -693 -29 -659
rect 29 -693 45 -659
rect 1613 -693 1629 -659
rect 1687 -693 1703 -659
rect 3271 -693 3287 -659
rect 3345 -693 3361 -659
rect 4929 -693 4945 -659
rect -5125 -797 -5091 -735
rect 5091 -797 5125 -735
rect -5125 -831 -5029 -797
rect 5029 -831 5125 -797
<< viali >>
rect -4991 495 -4957 671
rect -3333 495 -3299 671
rect -1675 495 -1641 671
rect -17 495 17 671
rect 1641 495 1675 671
rect 3299 495 3333 671
rect 4957 495 4991 671
rect -4929 402 -3361 436
rect -3271 402 -1703 436
rect -1613 402 -45 436
rect 45 402 1613 436
rect 1703 402 3271 436
rect 3361 402 4929 436
rect -4991 130 -4957 306
rect -3333 130 -3299 306
rect -1675 130 -1641 306
rect -17 130 17 306
rect 1641 130 1675 306
rect 3299 130 3333 306
rect 4957 130 4991 306
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect -4991 -235 -4957 -59
rect -3333 -235 -3299 -59
rect -1675 -235 -1641 -59
rect -17 -235 17 -59
rect 1641 -235 1675 -59
rect 3299 -235 3333 -59
rect 4957 -235 4991 -59
rect -4929 -328 -3361 -294
rect -3271 -328 -1703 -294
rect -1613 -328 -45 -294
rect 45 -328 1613 -294
rect 1703 -328 3271 -294
rect 3361 -328 4929 -294
rect -4991 -600 -4957 -424
rect -3333 -600 -3299 -424
rect -1675 -600 -1641 -424
rect -17 -600 17 -424
rect 1641 -600 1675 -424
rect 3299 -600 3333 -424
rect 4957 -600 4991 -424
rect -4929 -693 -3361 -659
rect -3271 -693 -1703 -659
rect -1613 -693 -45 -659
rect 45 -693 1613 -659
rect 1703 -693 3271 -659
rect 3361 -693 4929 -659
<< metal1 >>
rect -4997 671 -4951 683
rect -4997 495 -4991 671
rect -4957 495 -4951 671
rect -4997 483 -4951 495
rect -3339 671 -3293 683
rect -3339 495 -3333 671
rect -3299 495 -3293 671
rect -3339 483 -3293 495
rect -1681 671 -1635 683
rect -1681 495 -1675 671
rect -1641 495 -1635 671
rect -1681 483 -1635 495
rect -23 671 23 683
rect -23 495 -17 671
rect 17 495 23 671
rect -23 483 23 495
rect 1635 671 1681 683
rect 1635 495 1641 671
rect 1675 495 1681 671
rect 1635 483 1681 495
rect 3293 671 3339 683
rect 3293 495 3299 671
rect 3333 495 3339 671
rect 3293 483 3339 495
rect 4951 671 4997 683
rect 4951 495 4957 671
rect 4991 495 4997 671
rect 4951 483 4997 495
rect -4941 436 -3349 442
rect -4941 402 -4929 436
rect -3361 402 -3349 436
rect -4941 396 -3349 402
rect -3283 436 -1691 442
rect -3283 402 -3271 436
rect -1703 402 -1691 436
rect -3283 396 -1691 402
rect -1625 436 -33 442
rect -1625 402 -1613 436
rect -45 402 -33 436
rect -1625 396 -33 402
rect 33 436 1625 442
rect 33 402 45 436
rect 1613 402 1625 436
rect 33 396 1625 402
rect 1691 436 3283 442
rect 1691 402 1703 436
rect 3271 402 3283 436
rect 1691 396 3283 402
rect 3349 436 4941 442
rect 3349 402 3361 436
rect 4929 402 4941 436
rect 3349 396 4941 402
rect -4997 306 -4951 318
rect -4997 130 -4991 306
rect -4957 130 -4951 306
rect -4997 118 -4951 130
rect -3339 306 -3293 318
rect -3339 130 -3333 306
rect -3299 130 -3293 306
rect -3339 118 -3293 130
rect -1681 306 -1635 318
rect -1681 130 -1675 306
rect -1641 130 -1635 306
rect -1681 118 -1635 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 1635 306 1681 318
rect 1635 130 1641 306
rect 1675 130 1681 306
rect 1635 118 1681 130
rect 3293 306 3339 318
rect 3293 130 3299 306
rect 3333 130 3339 306
rect 3293 118 3339 130
rect 4951 306 4997 318
rect 4951 130 4957 306
rect 4991 130 4997 306
rect 4951 118 4997 130
rect -4941 71 -3349 77
rect -4941 37 -4929 71
rect -3361 37 -3349 71
rect -4941 31 -3349 37
rect -3283 71 -1691 77
rect -3283 37 -3271 71
rect -1703 37 -1691 71
rect -3283 31 -1691 37
rect -1625 71 -33 77
rect -1625 37 -1613 71
rect -45 37 -33 71
rect -1625 31 -33 37
rect 33 71 1625 77
rect 33 37 45 71
rect 1613 37 1625 71
rect 33 31 1625 37
rect 1691 71 3283 77
rect 1691 37 1703 71
rect 3271 37 3283 71
rect 1691 31 3283 37
rect 3349 71 4941 77
rect 3349 37 3361 71
rect 4929 37 4941 71
rect 3349 31 4941 37
rect -4997 -59 -4951 -47
rect -4997 -235 -4991 -59
rect -4957 -235 -4951 -59
rect -4997 -247 -4951 -235
rect -3339 -59 -3293 -47
rect -3339 -235 -3333 -59
rect -3299 -235 -3293 -59
rect -3339 -247 -3293 -235
rect -1681 -59 -1635 -47
rect -1681 -235 -1675 -59
rect -1641 -235 -1635 -59
rect -1681 -247 -1635 -235
rect -23 -59 23 -47
rect -23 -235 -17 -59
rect 17 -235 23 -59
rect -23 -247 23 -235
rect 1635 -59 1681 -47
rect 1635 -235 1641 -59
rect 1675 -235 1681 -59
rect 1635 -247 1681 -235
rect 3293 -59 3339 -47
rect 3293 -235 3299 -59
rect 3333 -235 3339 -59
rect 3293 -247 3339 -235
rect 4951 -59 4997 -47
rect 4951 -235 4957 -59
rect 4991 -235 4997 -59
rect 4951 -247 4997 -235
rect -4941 -294 -3349 -288
rect -4941 -328 -4929 -294
rect -3361 -328 -3349 -294
rect -4941 -334 -3349 -328
rect -3283 -294 -1691 -288
rect -3283 -328 -3271 -294
rect -1703 -328 -1691 -294
rect -3283 -334 -1691 -328
rect -1625 -294 -33 -288
rect -1625 -328 -1613 -294
rect -45 -328 -33 -294
rect -1625 -334 -33 -328
rect 33 -294 1625 -288
rect 33 -328 45 -294
rect 1613 -328 1625 -294
rect 33 -334 1625 -328
rect 1691 -294 3283 -288
rect 1691 -328 1703 -294
rect 3271 -328 3283 -294
rect 1691 -334 3283 -328
rect 3349 -294 4941 -288
rect 3349 -328 3361 -294
rect 4929 -328 4941 -294
rect 3349 -334 4941 -328
rect -4997 -424 -4951 -412
rect -4997 -600 -4991 -424
rect -4957 -600 -4951 -424
rect -4997 -612 -4951 -600
rect -3339 -424 -3293 -412
rect -3339 -600 -3333 -424
rect -3299 -600 -3293 -424
rect -3339 -612 -3293 -600
rect -1681 -424 -1635 -412
rect -1681 -600 -1675 -424
rect -1641 -600 -1635 -424
rect -1681 -612 -1635 -600
rect -23 -424 23 -412
rect -23 -600 -17 -424
rect 17 -600 23 -424
rect -23 -612 23 -600
rect 1635 -424 1681 -412
rect 1635 -600 1641 -424
rect 1675 -600 1681 -424
rect 1635 -612 1681 -600
rect 3293 -424 3339 -412
rect 3293 -600 3299 -424
rect 3333 -600 3339 -424
rect 3293 -612 3339 -600
rect 4951 -424 4997 -412
rect 4951 -600 4957 -424
rect 4991 -600 4997 -424
rect 4951 -612 4997 -600
rect -4941 -659 -3349 -653
rect -4941 -693 -4929 -659
rect -3361 -693 -3349 -659
rect -4941 -699 -3349 -693
rect -3283 -659 -1691 -653
rect -3283 -693 -3271 -659
rect -1703 -693 -1691 -659
rect -3283 -699 -1691 -693
rect -1625 -659 -33 -653
rect -1625 -693 -1613 -659
rect -45 -693 -33 -659
rect -1625 -699 -33 -693
rect 33 -659 1625 -653
rect 33 -693 45 -659
rect 1613 -693 1625 -659
rect 33 -699 1625 -693
rect 1691 -659 3283 -653
rect 1691 -693 1703 -659
rect 3271 -693 3283 -659
rect 1691 -699 3283 -693
rect 3349 -659 4941 -653
rect 3349 -693 3361 -659
rect 4929 -693 4941 -659
rect 3349 -699 4941 -693
<< properties >>
string FIXED_BBOX -5108 -814 5108 814
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 8 m 4 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712467038
<< nwell >>
rect -4412 -762 4412 762
<< mvpmos >>
rect -4154 -536 -4034 464
rect -3976 -536 -3856 464
rect -3798 -536 -3678 464
rect -3620 -536 -3500 464
rect -3442 -536 -3322 464
rect -3264 -536 -3144 464
rect -3086 -536 -2966 464
rect -2908 -536 -2788 464
rect -2730 -536 -2610 464
rect -2552 -536 -2432 464
rect -2374 -536 -2254 464
rect -2196 -536 -2076 464
rect -2018 -536 -1898 464
rect -1840 -536 -1720 464
rect -1662 -536 -1542 464
rect -1484 -536 -1364 464
rect -1306 -536 -1186 464
rect -1128 -536 -1008 464
rect -950 -536 -830 464
rect -772 -536 -652 464
rect -594 -536 -474 464
rect -416 -536 -296 464
rect -238 -536 -118 464
rect -60 -536 60 464
rect 118 -536 238 464
rect 296 -536 416 464
rect 474 -536 594 464
rect 652 -536 772 464
rect 830 -536 950 464
rect 1008 -536 1128 464
rect 1186 -536 1306 464
rect 1364 -536 1484 464
rect 1542 -536 1662 464
rect 1720 -536 1840 464
rect 1898 -536 2018 464
rect 2076 -536 2196 464
rect 2254 -536 2374 464
rect 2432 -536 2552 464
rect 2610 -536 2730 464
rect 2788 -536 2908 464
rect 2966 -536 3086 464
rect 3144 -536 3264 464
rect 3322 -536 3442 464
rect 3500 -536 3620 464
rect 3678 -536 3798 464
rect 3856 -536 3976 464
rect 4034 -536 4154 464
<< mvpdiff >>
rect -4212 452 -4154 464
rect -4212 -524 -4200 452
rect -4166 -524 -4154 452
rect -4212 -536 -4154 -524
rect -4034 452 -3976 464
rect -4034 -524 -4022 452
rect -3988 -524 -3976 452
rect -4034 -536 -3976 -524
rect -3856 452 -3798 464
rect -3856 -524 -3844 452
rect -3810 -524 -3798 452
rect -3856 -536 -3798 -524
rect -3678 452 -3620 464
rect -3678 -524 -3666 452
rect -3632 -524 -3620 452
rect -3678 -536 -3620 -524
rect -3500 452 -3442 464
rect -3500 -524 -3488 452
rect -3454 -524 -3442 452
rect -3500 -536 -3442 -524
rect -3322 452 -3264 464
rect -3322 -524 -3310 452
rect -3276 -524 -3264 452
rect -3322 -536 -3264 -524
rect -3144 452 -3086 464
rect -3144 -524 -3132 452
rect -3098 -524 -3086 452
rect -3144 -536 -3086 -524
rect -2966 452 -2908 464
rect -2966 -524 -2954 452
rect -2920 -524 -2908 452
rect -2966 -536 -2908 -524
rect -2788 452 -2730 464
rect -2788 -524 -2776 452
rect -2742 -524 -2730 452
rect -2788 -536 -2730 -524
rect -2610 452 -2552 464
rect -2610 -524 -2598 452
rect -2564 -524 -2552 452
rect -2610 -536 -2552 -524
rect -2432 452 -2374 464
rect -2432 -524 -2420 452
rect -2386 -524 -2374 452
rect -2432 -536 -2374 -524
rect -2254 452 -2196 464
rect -2254 -524 -2242 452
rect -2208 -524 -2196 452
rect -2254 -536 -2196 -524
rect -2076 452 -2018 464
rect -2076 -524 -2064 452
rect -2030 -524 -2018 452
rect -2076 -536 -2018 -524
rect -1898 452 -1840 464
rect -1898 -524 -1886 452
rect -1852 -524 -1840 452
rect -1898 -536 -1840 -524
rect -1720 452 -1662 464
rect -1720 -524 -1708 452
rect -1674 -524 -1662 452
rect -1720 -536 -1662 -524
rect -1542 452 -1484 464
rect -1542 -524 -1530 452
rect -1496 -524 -1484 452
rect -1542 -536 -1484 -524
rect -1364 452 -1306 464
rect -1364 -524 -1352 452
rect -1318 -524 -1306 452
rect -1364 -536 -1306 -524
rect -1186 452 -1128 464
rect -1186 -524 -1174 452
rect -1140 -524 -1128 452
rect -1186 -536 -1128 -524
rect -1008 452 -950 464
rect -1008 -524 -996 452
rect -962 -524 -950 452
rect -1008 -536 -950 -524
rect -830 452 -772 464
rect -830 -524 -818 452
rect -784 -524 -772 452
rect -830 -536 -772 -524
rect -652 452 -594 464
rect -652 -524 -640 452
rect -606 -524 -594 452
rect -652 -536 -594 -524
rect -474 452 -416 464
rect -474 -524 -462 452
rect -428 -524 -416 452
rect -474 -536 -416 -524
rect -296 452 -238 464
rect -296 -524 -284 452
rect -250 -524 -238 452
rect -296 -536 -238 -524
rect -118 452 -60 464
rect -118 -524 -106 452
rect -72 -524 -60 452
rect -118 -536 -60 -524
rect 60 452 118 464
rect 60 -524 72 452
rect 106 -524 118 452
rect 60 -536 118 -524
rect 238 452 296 464
rect 238 -524 250 452
rect 284 -524 296 452
rect 238 -536 296 -524
rect 416 452 474 464
rect 416 -524 428 452
rect 462 -524 474 452
rect 416 -536 474 -524
rect 594 452 652 464
rect 594 -524 606 452
rect 640 -524 652 452
rect 594 -536 652 -524
rect 772 452 830 464
rect 772 -524 784 452
rect 818 -524 830 452
rect 772 -536 830 -524
rect 950 452 1008 464
rect 950 -524 962 452
rect 996 -524 1008 452
rect 950 -536 1008 -524
rect 1128 452 1186 464
rect 1128 -524 1140 452
rect 1174 -524 1186 452
rect 1128 -536 1186 -524
rect 1306 452 1364 464
rect 1306 -524 1318 452
rect 1352 -524 1364 452
rect 1306 -536 1364 -524
rect 1484 452 1542 464
rect 1484 -524 1496 452
rect 1530 -524 1542 452
rect 1484 -536 1542 -524
rect 1662 452 1720 464
rect 1662 -524 1674 452
rect 1708 -524 1720 452
rect 1662 -536 1720 -524
rect 1840 452 1898 464
rect 1840 -524 1852 452
rect 1886 -524 1898 452
rect 1840 -536 1898 -524
rect 2018 452 2076 464
rect 2018 -524 2030 452
rect 2064 -524 2076 452
rect 2018 -536 2076 -524
rect 2196 452 2254 464
rect 2196 -524 2208 452
rect 2242 -524 2254 452
rect 2196 -536 2254 -524
rect 2374 452 2432 464
rect 2374 -524 2386 452
rect 2420 -524 2432 452
rect 2374 -536 2432 -524
rect 2552 452 2610 464
rect 2552 -524 2564 452
rect 2598 -524 2610 452
rect 2552 -536 2610 -524
rect 2730 452 2788 464
rect 2730 -524 2742 452
rect 2776 -524 2788 452
rect 2730 -536 2788 -524
rect 2908 452 2966 464
rect 2908 -524 2920 452
rect 2954 -524 2966 452
rect 2908 -536 2966 -524
rect 3086 452 3144 464
rect 3086 -524 3098 452
rect 3132 -524 3144 452
rect 3086 -536 3144 -524
rect 3264 452 3322 464
rect 3264 -524 3276 452
rect 3310 -524 3322 452
rect 3264 -536 3322 -524
rect 3442 452 3500 464
rect 3442 -524 3454 452
rect 3488 -524 3500 452
rect 3442 -536 3500 -524
rect 3620 452 3678 464
rect 3620 -524 3632 452
rect 3666 -524 3678 452
rect 3620 -536 3678 -524
rect 3798 452 3856 464
rect 3798 -524 3810 452
rect 3844 -524 3856 452
rect 3798 -536 3856 -524
rect 3976 452 4034 464
rect 3976 -524 3988 452
rect 4022 -524 4034 452
rect 3976 -536 4034 -524
rect 4154 452 4212 464
rect 4154 -524 4166 452
rect 4200 -524 4212 452
rect 4154 -536 4212 -524
<< mvpdiffc >>
rect -4200 -524 -4166 452
rect -4022 -524 -3988 452
rect -3844 -524 -3810 452
rect -3666 -524 -3632 452
rect -3488 -524 -3454 452
rect -3310 -524 -3276 452
rect -3132 -524 -3098 452
rect -2954 -524 -2920 452
rect -2776 -524 -2742 452
rect -2598 -524 -2564 452
rect -2420 -524 -2386 452
rect -2242 -524 -2208 452
rect -2064 -524 -2030 452
rect -1886 -524 -1852 452
rect -1708 -524 -1674 452
rect -1530 -524 -1496 452
rect -1352 -524 -1318 452
rect -1174 -524 -1140 452
rect -996 -524 -962 452
rect -818 -524 -784 452
rect -640 -524 -606 452
rect -462 -524 -428 452
rect -284 -524 -250 452
rect -106 -524 -72 452
rect 72 -524 106 452
rect 250 -524 284 452
rect 428 -524 462 452
rect 606 -524 640 452
rect 784 -524 818 452
rect 962 -524 996 452
rect 1140 -524 1174 452
rect 1318 -524 1352 452
rect 1496 -524 1530 452
rect 1674 -524 1708 452
rect 1852 -524 1886 452
rect 2030 -524 2064 452
rect 2208 -524 2242 452
rect 2386 -524 2420 452
rect 2564 -524 2598 452
rect 2742 -524 2776 452
rect 2920 -524 2954 452
rect 3098 -524 3132 452
rect 3276 -524 3310 452
rect 3454 -524 3488 452
rect 3632 -524 3666 452
rect 3810 -524 3844 452
rect 3988 -524 4022 452
rect 4166 -524 4200 452
<< mvnsubdiff >>
rect -4346 684 4346 696
rect -4346 650 -4238 684
rect 4238 650 4346 684
rect -4346 638 4346 650
rect -4346 588 -4288 638
rect -4346 -588 -4334 588
rect -4300 -588 -4288 588
rect 4288 588 4346 638
rect -4346 -638 -4288 -588
rect 4288 -588 4300 588
rect 4334 -588 4346 588
rect 4288 -638 4346 -588
rect -4346 -650 4346 -638
rect -4346 -684 -4238 -650
rect 4238 -684 4346 -650
rect -4346 -696 4346 -684
<< mvnsubdiffcont >>
rect -4238 650 4238 684
rect -4334 -588 -4300 588
rect 4300 -588 4334 588
rect -4238 -684 4238 -650
<< poly >>
rect -4154 545 -4034 561
rect -4154 511 -4138 545
rect -4050 511 -4034 545
rect -4154 464 -4034 511
rect -3976 545 -3856 561
rect -3976 511 -3960 545
rect -3872 511 -3856 545
rect -3976 464 -3856 511
rect -3798 545 -3678 561
rect -3798 511 -3782 545
rect -3694 511 -3678 545
rect -3798 464 -3678 511
rect -3620 545 -3500 561
rect -3620 511 -3604 545
rect -3516 511 -3500 545
rect -3620 464 -3500 511
rect -3442 545 -3322 561
rect -3442 511 -3426 545
rect -3338 511 -3322 545
rect -3442 464 -3322 511
rect -3264 545 -3144 561
rect -3264 511 -3248 545
rect -3160 511 -3144 545
rect -3264 464 -3144 511
rect -3086 545 -2966 561
rect -3086 511 -3070 545
rect -2982 511 -2966 545
rect -3086 464 -2966 511
rect -2908 545 -2788 561
rect -2908 511 -2892 545
rect -2804 511 -2788 545
rect -2908 464 -2788 511
rect -2730 545 -2610 561
rect -2730 511 -2714 545
rect -2626 511 -2610 545
rect -2730 464 -2610 511
rect -2552 545 -2432 561
rect -2552 511 -2536 545
rect -2448 511 -2432 545
rect -2552 464 -2432 511
rect -2374 545 -2254 561
rect -2374 511 -2358 545
rect -2270 511 -2254 545
rect -2374 464 -2254 511
rect -2196 545 -2076 561
rect -2196 511 -2180 545
rect -2092 511 -2076 545
rect -2196 464 -2076 511
rect -2018 545 -1898 561
rect -2018 511 -2002 545
rect -1914 511 -1898 545
rect -2018 464 -1898 511
rect -1840 545 -1720 561
rect -1840 511 -1824 545
rect -1736 511 -1720 545
rect -1840 464 -1720 511
rect -1662 545 -1542 561
rect -1662 511 -1646 545
rect -1558 511 -1542 545
rect -1662 464 -1542 511
rect -1484 545 -1364 561
rect -1484 511 -1468 545
rect -1380 511 -1364 545
rect -1484 464 -1364 511
rect -1306 545 -1186 561
rect -1306 511 -1290 545
rect -1202 511 -1186 545
rect -1306 464 -1186 511
rect -1128 545 -1008 561
rect -1128 511 -1112 545
rect -1024 511 -1008 545
rect -1128 464 -1008 511
rect -950 545 -830 561
rect -950 511 -934 545
rect -846 511 -830 545
rect -950 464 -830 511
rect -772 545 -652 561
rect -772 511 -756 545
rect -668 511 -652 545
rect -772 464 -652 511
rect -594 545 -474 561
rect -594 511 -578 545
rect -490 511 -474 545
rect -594 464 -474 511
rect -416 545 -296 561
rect -416 511 -400 545
rect -312 511 -296 545
rect -416 464 -296 511
rect -238 545 -118 561
rect -238 511 -222 545
rect -134 511 -118 545
rect -238 464 -118 511
rect -60 545 60 561
rect -60 511 -44 545
rect 44 511 60 545
rect -60 464 60 511
rect 118 545 238 561
rect 118 511 134 545
rect 222 511 238 545
rect 118 464 238 511
rect 296 545 416 561
rect 296 511 312 545
rect 400 511 416 545
rect 296 464 416 511
rect 474 545 594 561
rect 474 511 490 545
rect 578 511 594 545
rect 474 464 594 511
rect 652 545 772 561
rect 652 511 668 545
rect 756 511 772 545
rect 652 464 772 511
rect 830 545 950 561
rect 830 511 846 545
rect 934 511 950 545
rect 830 464 950 511
rect 1008 545 1128 561
rect 1008 511 1024 545
rect 1112 511 1128 545
rect 1008 464 1128 511
rect 1186 545 1306 561
rect 1186 511 1202 545
rect 1290 511 1306 545
rect 1186 464 1306 511
rect 1364 545 1484 561
rect 1364 511 1380 545
rect 1468 511 1484 545
rect 1364 464 1484 511
rect 1542 545 1662 561
rect 1542 511 1558 545
rect 1646 511 1662 545
rect 1542 464 1662 511
rect 1720 545 1840 561
rect 1720 511 1736 545
rect 1824 511 1840 545
rect 1720 464 1840 511
rect 1898 545 2018 561
rect 1898 511 1914 545
rect 2002 511 2018 545
rect 1898 464 2018 511
rect 2076 545 2196 561
rect 2076 511 2092 545
rect 2180 511 2196 545
rect 2076 464 2196 511
rect 2254 545 2374 561
rect 2254 511 2270 545
rect 2358 511 2374 545
rect 2254 464 2374 511
rect 2432 545 2552 561
rect 2432 511 2448 545
rect 2536 511 2552 545
rect 2432 464 2552 511
rect 2610 545 2730 561
rect 2610 511 2626 545
rect 2714 511 2730 545
rect 2610 464 2730 511
rect 2788 545 2908 561
rect 2788 511 2804 545
rect 2892 511 2908 545
rect 2788 464 2908 511
rect 2966 545 3086 561
rect 2966 511 2982 545
rect 3070 511 3086 545
rect 2966 464 3086 511
rect 3144 545 3264 561
rect 3144 511 3160 545
rect 3248 511 3264 545
rect 3144 464 3264 511
rect 3322 545 3442 561
rect 3322 511 3338 545
rect 3426 511 3442 545
rect 3322 464 3442 511
rect 3500 545 3620 561
rect 3500 511 3516 545
rect 3604 511 3620 545
rect 3500 464 3620 511
rect 3678 545 3798 561
rect 3678 511 3694 545
rect 3782 511 3798 545
rect 3678 464 3798 511
rect 3856 545 3976 561
rect 3856 511 3872 545
rect 3960 511 3976 545
rect 3856 464 3976 511
rect 4034 545 4154 561
rect 4034 511 4050 545
rect 4138 511 4154 545
rect 4034 464 4154 511
rect -4154 -562 -4034 -536
rect -3976 -562 -3856 -536
rect -3798 -562 -3678 -536
rect -3620 -562 -3500 -536
rect -3442 -562 -3322 -536
rect -3264 -562 -3144 -536
rect -3086 -562 -2966 -536
rect -2908 -562 -2788 -536
rect -2730 -562 -2610 -536
rect -2552 -562 -2432 -536
rect -2374 -562 -2254 -536
rect -2196 -562 -2076 -536
rect -2018 -562 -1898 -536
rect -1840 -562 -1720 -536
rect -1662 -562 -1542 -536
rect -1484 -562 -1364 -536
rect -1306 -562 -1186 -536
rect -1128 -562 -1008 -536
rect -950 -562 -830 -536
rect -772 -562 -652 -536
rect -594 -562 -474 -536
rect -416 -562 -296 -536
rect -238 -562 -118 -536
rect -60 -562 60 -536
rect 118 -562 238 -536
rect 296 -562 416 -536
rect 474 -562 594 -536
rect 652 -562 772 -536
rect 830 -562 950 -536
rect 1008 -562 1128 -536
rect 1186 -562 1306 -536
rect 1364 -562 1484 -536
rect 1542 -562 1662 -536
rect 1720 -562 1840 -536
rect 1898 -562 2018 -536
rect 2076 -562 2196 -536
rect 2254 -562 2374 -536
rect 2432 -562 2552 -536
rect 2610 -562 2730 -536
rect 2788 -562 2908 -536
rect 2966 -562 3086 -536
rect 3144 -562 3264 -536
rect 3322 -562 3442 -536
rect 3500 -562 3620 -536
rect 3678 -562 3798 -536
rect 3856 -562 3976 -536
rect 4034 -562 4154 -536
<< polycont >>
rect -4138 511 -4050 545
rect -3960 511 -3872 545
rect -3782 511 -3694 545
rect -3604 511 -3516 545
rect -3426 511 -3338 545
rect -3248 511 -3160 545
rect -3070 511 -2982 545
rect -2892 511 -2804 545
rect -2714 511 -2626 545
rect -2536 511 -2448 545
rect -2358 511 -2270 545
rect -2180 511 -2092 545
rect -2002 511 -1914 545
rect -1824 511 -1736 545
rect -1646 511 -1558 545
rect -1468 511 -1380 545
rect -1290 511 -1202 545
rect -1112 511 -1024 545
rect -934 511 -846 545
rect -756 511 -668 545
rect -578 511 -490 545
rect -400 511 -312 545
rect -222 511 -134 545
rect -44 511 44 545
rect 134 511 222 545
rect 312 511 400 545
rect 490 511 578 545
rect 668 511 756 545
rect 846 511 934 545
rect 1024 511 1112 545
rect 1202 511 1290 545
rect 1380 511 1468 545
rect 1558 511 1646 545
rect 1736 511 1824 545
rect 1914 511 2002 545
rect 2092 511 2180 545
rect 2270 511 2358 545
rect 2448 511 2536 545
rect 2626 511 2714 545
rect 2804 511 2892 545
rect 2982 511 3070 545
rect 3160 511 3248 545
rect 3338 511 3426 545
rect 3516 511 3604 545
rect 3694 511 3782 545
rect 3872 511 3960 545
rect 4050 511 4138 545
<< locali >>
rect -4334 650 -4238 684
rect 4238 650 4334 684
rect -4334 588 -4300 650
rect 4300 588 4334 650
rect -4154 511 -4138 545
rect -4050 511 -4034 545
rect -3976 511 -3960 545
rect -3872 511 -3856 545
rect -3798 511 -3782 545
rect -3694 511 -3678 545
rect -3620 511 -3604 545
rect -3516 511 -3500 545
rect -3442 511 -3426 545
rect -3338 511 -3322 545
rect -3264 511 -3248 545
rect -3160 511 -3144 545
rect -3086 511 -3070 545
rect -2982 511 -2966 545
rect -2908 511 -2892 545
rect -2804 511 -2788 545
rect -2730 511 -2714 545
rect -2626 511 -2610 545
rect -2552 511 -2536 545
rect -2448 511 -2432 545
rect -2374 511 -2358 545
rect -2270 511 -2254 545
rect -2196 511 -2180 545
rect -2092 511 -2076 545
rect -2018 511 -2002 545
rect -1914 511 -1898 545
rect -1840 511 -1824 545
rect -1736 511 -1720 545
rect -1662 511 -1646 545
rect -1558 511 -1542 545
rect -1484 511 -1468 545
rect -1380 511 -1364 545
rect -1306 511 -1290 545
rect -1202 511 -1186 545
rect -1128 511 -1112 545
rect -1024 511 -1008 545
rect -950 511 -934 545
rect -846 511 -830 545
rect -772 511 -756 545
rect -668 511 -652 545
rect -594 511 -578 545
rect -490 511 -474 545
rect -416 511 -400 545
rect -312 511 -296 545
rect -238 511 -222 545
rect -134 511 -118 545
rect -60 511 -44 545
rect 44 511 60 545
rect 118 511 134 545
rect 222 511 238 545
rect 296 511 312 545
rect 400 511 416 545
rect 474 511 490 545
rect 578 511 594 545
rect 652 511 668 545
rect 756 511 772 545
rect 830 511 846 545
rect 934 511 950 545
rect 1008 511 1024 545
rect 1112 511 1128 545
rect 1186 511 1202 545
rect 1290 511 1306 545
rect 1364 511 1380 545
rect 1468 511 1484 545
rect 1542 511 1558 545
rect 1646 511 1662 545
rect 1720 511 1736 545
rect 1824 511 1840 545
rect 1898 511 1914 545
rect 2002 511 2018 545
rect 2076 511 2092 545
rect 2180 511 2196 545
rect 2254 511 2270 545
rect 2358 511 2374 545
rect 2432 511 2448 545
rect 2536 511 2552 545
rect 2610 511 2626 545
rect 2714 511 2730 545
rect 2788 511 2804 545
rect 2892 511 2908 545
rect 2966 511 2982 545
rect 3070 511 3086 545
rect 3144 511 3160 545
rect 3248 511 3264 545
rect 3322 511 3338 545
rect 3426 511 3442 545
rect 3500 511 3516 545
rect 3604 511 3620 545
rect 3678 511 3694 545
rect 3782 511 3798 545
rect 3856 511 3872 545
rect 3960 511 3976 545
rect 4034 511 4050 545
rect 4138 511 4154 545
rect -4200 452 -4166 468
rect -4200 -540 -4166 -524
rect -4022 452 -3988 468
rect -4022 -540 -3988 -524
rect -3844 452 -3810 468
rect -3844 -540 -3810 -524
rect -3666 452 -3632 468
rect -3666 -540 -3632 -524
rect -3488 452 -3454 468
rect -3488 -540 -3454 -524
rect -3310 452 -3276 468
rect -3310 -540 -3276 -524
rect -3132 452 -3098 468
rect -3132 -540 -3098 -524
rect -2954 452 -2920 468
rect -2954 -540 -2920 -524
rect -2776 452 -2742 468
rect -2776 -540 -2742 -524
rect -2598 452 -2564 468
rect -2598 -540 -2564 -524
rect -2420 452 -2386 468
rect -2420 -540 -2386 -524
rect -2242 452 -2208 468
rect -2242 -540 -2208 -524
rect -2064 452 -2030 468
rect -2064 -540 -2030 -524
rect -1886 452 -1852 468
rect -1886 -540 -1852 -524
rect -1708 452 -1674 468
rect -1708 -540 -1674 -524
rect -1530 452 -1496 468
rect -1530 -540 -1496 -524
rect -1352 452 -1318 468
rect -1352 -540 -1318 -524
rect -1174 452 -1140 468
rect -1174 -540 -1140 -524
rect -996 452 -962 468
rect -996 -540 -962 -524
rect -818 452 -784 468
rect -818 -540 -784 -524
rect -640 452 -606 468
rect -640 -540 -606 -524
rect -462 452 -428 468
rect -462 -540 -428 -524
rect -284 452 -250 468
rect -284 -540 -250 -524
rect -106 452 -72 468
rect -106 -540 -72 -524
rect 72 452 106 468
rect 72 -540 106 -524
rect 250 452 284 468
rect 250 -540 284 -524
rect 428 452 462 468
rect 428 -540 462 -524
rect 606 452 640 468
rect 606 -540 640 -524
rect 784 452 818 468
rect 784 -540 818 -524
rect 962 452 996 468
rect 962 -540 996 -524
rect 1140 452 1174 468
rect 1140 -540 1174 -524
rect 1318 452 1352 468
rect 1318 -540 1352 -524
rect 1496 452 1530 468
rect 1496 -540 1530 -524
rect 1674 452 1708 468
rect 1674 -540 1708 -524
rect 1852 452 1886 468
rect 1852 -540 1886 -524
rect 2030 452 2064 468
rect 2030 -540 2064 -524
rect 2208 452 2242 468
rect 2208 -540 2242 -524
rect 2386 452 2420 468
rect 2386 -540 2420 -524
rect 2564 452 2598 468
rect 2564 -540 2598 -524
rect 2742 452 2776 468
rect 2742 -540 2776 -524
rect 2920 452 2954 468
rect 2920 -540 2954 -524
rect 3098 452 3132 468
rect 3098 -540 3132 -524
rect 3276 452 3310 468
rect 3276 -540 3310 -524
rect 3454 452 3488 468
rect 3454 -540 3488 -524
rect 3632 452 3666 468
rect 3632 -540 3666 -524
rect 3810 452 3844 468
rect 3810 -540 3844 -524
rect 3988 452 4022 468
rect 3988 -540 4022 -524
rect 4166 452 4200 468
rect 4166 -540 4200 -524
rect -4334 -650 -4300 -588
rect 4300 -650 4334 -588
rect -4334 -684 -4238 -650
rect 4238 -684 4334 -650
<< viali >>
rect -4138 511 -4050 545
rect -3960 511 -3872 545
rect -3782 511 -3694 545
rect -3604 511 -3516 545
rect -3426 511 -3338 545
rect -3248 511 -3160 545
rect -3070 511 -2982 545
rect -2892 511 -2804 545
rect -2714 511 -2626 545
rect -2536 511 -2448 545
rect -2358 511 -2270 545
rect -2180 511 -2092 545
rect -2002 511 -1914 545
rect -1824 511 -1736 545
rect -1646 511 -1558 545
rect -1468 511 -1380 545
rect -1290 511 -1202 545
rect -1112 511 -1024 545
rect -934 511 -846 545
rect -756 511 -668 545
rect -578 511 -490 545
rect -400 511 -312 545
rect -222 511 -134 545
rect -44 511 44 545
rect 134 511 222 545
rect 312 511 400 545
rect 490 511 578 545
rect 668 511 756 545
rect 846 511 934 545
rect 1024 511 1112 545
rect 1202 511 1290 545
rect 1380 511 1468 545
rect 1558 511 1646 545
rect 1736 511 1824 545
rect 1914 511 2002 545
rect 2092 511 2180 545
rect 2270 511 2358 545
rect 2448 511 2536 545
rect 2626 511 2714 545
rect 2804 511 2892 545
rect 2982 511 3070 545
rect 3160 511 3248 545
rect 3338 511 3426 545
rect 3516 511 3604 545
rect 3694 511 3782 545
rect 3872 511 3960 545
rect 4050 511 4138 545
rect -4200 -524 -4166 452
rect -4022 -524 -3988 452
rect -3844 -524 -3810 452
rect -3666 -524 -3632 452
rect -3488 -524 -3454 452
rect -3310 -524 -3276 452
rect -3132 -524 -3098 452
rect -2954 -524 -2920 452
rect -2776 -524 -2742 452
rect -2598 -524 -2564 452
rect -2420 -524 -2386 452
rect -2242 -524 -2208 452
rect -2064 -524 -2030 452
rect -1886 -524 -1852 452
rect -1708 -524 -1674 452
rect -1530 -524 -1496 452
rect -1352 -524 -1318 452
rect -1174 -524 -1140 452
rect -996 -524 -962 452
rect -818 -524 -784 452
rect -640 -524 -606 452
rect -462 -524 -428 452
rect -284 -524 -250 452
rect -106 -524 -72 452
rect 72 -524 106 452
rect 250 -524 284 452
rect 428 -524 462 452
rect 606 -524 640 452
rect 784 -524 818 452
rect 962 -524 996 452
rect 1140 -524 1174 452
rect 1318 -524 1352 452
rect 1496 -524 1530 452
rect 1674 -524 1708 452
rect 1852 -524 1886 452
rect 2030 -524 2064 452
rect 2208 -524 2242 452
rect 2386 -524 2420 452
rect 2564 -524 2598 452
rect 2742 -524 2776 452
rect 2920 -524 2954 452
rect 3098 -524 3132 452
rect 3276 -524 3310 452
rect 3454 -524 3488 452
rect 3632 -524 3666 452
rect 3810 -524 3844 452
rect 3988 -524 4022 452
rect 4166 -524 4200 452
<< metal1 >>
rect -4150 545 -4038 551
rect -4150 511 -4138 545
rect -4050 511 -4038 545
rect -4150 505 -4038 511
rect -3972 545 -3860 551
rect -3972 511 -3960 545
rect -3872 511 -3860 545
rect -3972 505 -3860 511
rect -3794 545 -3682 551
rect -3794 511 -3782 545
rect -3694 511 -3682 545
rect -3794 505 -3682 511
rect -3616 545 -3504 551
rect -3616 511 -3604 545
rect -3516 511 -3504 545
rect -3616 505 -3504 511
rect -3438 545 -3326 551
rect -3438 511 -3426 545
rect -3338 511 -3326 545
rect -3438 505 -3326 511
rect -3260 545 -3148 551
rect -3260 511 -3248 545
rect -3160 511 -3148 545
rect -3260 505 -3148 511
rect -3082 545 -2970 551
rect -3082 511 -3070 545
rect -2982 511 -2970 545
rect -3082 505 -2970 511
rect -2904 545 -2792 551
rect -2904 511 -2892 545
rect -2804 511 -2792 545
rect -2904 505 -2792 511
rect -2726 545 -2614 551
rect -2726 511 -2714 545
rect -2626 511 -2614 545
rect -2726 505 -2614 511
rect -2548 545 -2436 551
rect -2548 511 -2536 545
rect -2448 511 -2436 545
rect -2548 505 -2436 511
rect -2370 545 -2258 551
rect -2370 511 -2358 545
rect -2270 511 -2258 545
rect -2370 505 -2258 511
rect -2192 545 -2080 551
rect -2192 511 -2180 545
rect -2092 511 -2080 545
rect -2192 505 -2080 511
rect -2014 545 -1902 551
rect -2014 511 -2002 545
rect -1914 511 -1902 545
rect -2014 505 -1902 511
rect -1836 545 -1724 551
rect -1836 511 -1824 545
rect -1736 511 -1724 545
rect -1836 505 -1724 511
rect -1658 545 -1546 551
rect -1658 511 -1646 545
rect -1558 511 -1546 545
rect -1658 505 -1546 511
rect -1480 545 -1368 551
rect -1480 511 -1468 545
rect -1380 511 -1368 545
rect -1480 505 -1368 511
rect -1302 545 -1190 551
rect -1302 511 -1290 545
rect -1202 511 -1190 545
rect -1302 505 -1190 511
rect -1124 545 -1012 551
rect -1124 511 -1112 545
rect -1024 511 -1012 545
rect -1124 505 -1012 511
rect -946 545 -834 551
rect -946 511 -934 545
rect -846 511 -834 545
rect -946 505 -834 511
rect -768 545 -656 551
rect -768 511 -756 545
rect -668 511 -656 545
rect -768 505 -656 511
rect -590 545 -478 551
rect -590 511 -578 545
rect -490 511 -478 545
rect -590 505 -478 511
rect -412 545 -300 551
rect -412 511 -400 545
rect -312 511 -300 545
rect -412 505 -300 511
rect -234 545 -122 551
rect -234 511 -222 545
rect -134 511 -122 545
rect -234 505 -122 511
rect -56 545 56 551
rect -56 511 -44 545
rect 44 511 56 545
rect -56 505 56 511
rect 122 545 234 551
rect 122 511 134 545
rect 222 511 234 545
rect 122 505 234 511
rect 300 545 412 551
rect 300 511 312 545
rect 400 511 412 545
rect 300 505 412 511
rect 478 545 590 551
rect 478 511 490 545
rect 578 511 590 545
rect 478 505 590 511
rect 656 545 768 551
rect 656 511 668 545
rect 756 511 768 545
rect 656 505 768 511
rect 834 545 946 551
rect 834 511 846 545
rect 934 511 946 545
rect 834 505 946 511
rect 1012 545 1124 551
rect 1012 511 1024 545
rect 1112 511 1124 545
rect 1012 505 1124 511
rect 1190 545 1302 551
rect 1190 511 1202 545
rect 1290 511 1302 545
rect 1190 505 1302 511
rect 1368 545 1480 551
rect 1368 511 1380 545
rect 1468 511 1480 545
rect 1368 505 1480 511
rect 1546 545 1658 551
rect 1546 511 1558 545
rect 1646 511 1658 545
rect 1546 505 1658 511
rect 1724 545 1836 551
rect 1724 511 1736 545
rect 1824 511 1836 545
rect 1724 505 1836 511
rect 1902 545 2014 551
rect 1902 511 1914 545
rect 2002 511 2014 545
rect 1902 505 2014 511
rect 2080 545 2192 551
rect 2080 511 2092 545
rect 2180 511 2192 545
rect 2080 505 2192 511
rect 2258 545 2370 551
rect 2258 511 2270 545
rect 2358 511 2370 545
rect 2258 505 2370 511
rect 2436 545 2548 551
rect 2436 511 2448 545
rect 2536 511 2548 545
rect 2436 505 2548 511
rect 2614 545 2726 551
rect 2614 511 2626 545
rect 2714 511 2726 545
rect 2614 505 2726 511
rect 2792 545 2904 551
rect 2792 511 2804 545
rect 2892 511 2904 545
rect 2792 505 2904 511
rect 2970 545 3082 551
rect 2970 511 2982 545
rect 3070 511 3082 545
rect 2970 505 3082 511
rect 3148 545 3260 551
rect 3148 511 3160 545
rect 3248 511 3260 545
rect 3148 505 3260 511
rect 3326 545 3438 551
rect 3326 511 3338 545
rect 3426 511 3438 545
rect 3326 505 3438 511
rect 3504 545 3616 551
rect 3504 511 3516 545
rect 3604 511 3616 545
rect 3504 505 3616 511
rect 3682 545 3794 551
rect 3682 511 3694 545
rect 3782 511 3794 545
rect 3682 505 3794 511
rect 3860 545 3972 551
rect 3860 511 3872 545
rect 3960 511 3972 545
rect 3860 505 3972 511
rect 4038 545 4150 551
rect 4038 511 4050 545
rect 4138 511 4150 545
rect 4038 505 4150 511
rect -4206 452 -4160 464
rect -4206 -524 -4200 452
rect -4166 -524 -4160 452
rect -4206 -536 -4160 -524
rect -4028 452 -3982 464
rect -4028 -524 -4022 452
rect -3988 -524 -3982 452
rect -4028 -536 -3982 -524
rect -3850 452 -3804 464
rect -3850 -524 -3844 452
rect -3810 -524 -3804 452
rect -3850 -536 -3804 -524
rect -3672 452 -3626 464
rect -3672 -524 -3666 452
rect -3632 -524 -3626 452
rect -3672 -536 -3626 -524
rect -3494 452 -3448 464
rect -3494 -524 -3488 452
rect -3454 -524 -3448 452
rect -3494 -536 -3448 -524
rect -3316 452 -3270 464
rect -3316 -524 -3310 452
rect -3276 -524 -3270 452
rect -3316 -536 -3270 -524
rect -3138 452 -3092 464
rect -3138 -524 -3132 452
rect -3098 -524 -3092 452
rect -3138 -536 -3092 -524
rect -2960 452 -2914 464
rect -2960 -524 -2954 452
rect -2920 -524 -2914 452
rect -2960 -536 -2914 -524
rect -2782 452 -2736 464
rect -2782 -524 -2776 452
rect -2742 -524 -2736 452
rect -2782 -536 -2736 -524
rect -2604 452 -2558 464
rect -2604 -524 -2598 452
rect -2564 -524 -2558 452
rect -2604 -536 -2558 -524
rect -2426 452 -2380 464
rect -2426 -524 -2420 452
rect -2386 -524 -2380 452
rect -2426 -536 -2380 -524
rect -2248 452 -2202 464
rect -2248 -524 -2242 452
rect -2208 -524 -2202 452
rect -2248 -536 -2202 -524
rect -2070 452 -2024 464
rect -2070 -524 -2064 452
rect -2030 -524 -2024 452
rect -2070 -536 -2024 -524
rect -1892 452 -1846 464
rect -1892 -524 -1886 452
rect -1852 -524 -1846 452
rect -1892 -536 -1846 -524
rect -1714 452 -1668 464
rect -1714 -524 -1708 452
rect -1674 -524 -1668 452
rect -1714 -536 -1668 -524
rect -1536 452 -1490 464
rect -1536 -524 -1530 452
rect -1496 -524 -1490 452
rect -1536 -536 -1490 -524
rect -1358 452 -1312 464
rect -1358 -524 -1352 452
rect -1318 -524 -1312 452
rect -1358 -536 -1312 -524
rect -1180 452 -1134 464
rect -1180 -524 -1174 452
rect -1140 -524 -1134 452
rect -1180 -536 -1134 -524
rect -1002 452 -956 464
rect -1002 -524 -996 452
rect -962 -524 -956 452
rect -1002 -536 -956 -524
rect -824 452 -778 464
rect -824 -524 -818 452
rect -784 -524 -778 452
rect -824 -536 -778 -524
rect -646 452 -600 464
rect -646 -524 -640 452
rect -606 -524 -600 452
rect -646 -536 -600 -524
rect -468 452 -422 464
rect -468 -524 -462 452
rect -428 -524 -422 452
rect -468 -536 -422 -524
rect -290 452 -244 464
rect -290 -524 -284 452
rect -250 -524 -244 452
rect -290 -536 -244 -524
rect -112 452 -66 464
rect -112 -524 -106 452
rect -72 -524 -66 452
rect -112 -536 -66 -524
rect 66 452 112 464
rect 66 -524 72 452
rect 106 -524 112 452
rect 66 -536 112 -524
rect 244 452 290 464
rect 244 -524 250 452
rect 284 -524 290 452
rect 244 -536 290 -524
rect 422 452 468 464
rect 422 -524 428 452
rect 462 -524 468 452
rect 422 -536 468 -524
rect 600 452 646 464
rect 600 -524 606 452
rect 640 -524 646 452
rect 600 -536 646 -524
rect 778 452 824 464
rect 778 -524 784 452
rect 818 -524 824 452
rect 778 -536 824 -524
rect 956 452 1002 464
rect 956 -524 962 452
rect 996 -524 1002 452
rect 956 -536 1002 -524
rect 1134 452 1180 464
rect 1134 -524 1140 452
rect 1174 -524 1180 452
rect 1134 -536 1180 -524
rect 1312 452 1358 464
rect 1312 -524 1318 452
rect 1352 -524 1358 452
rect 1312 -536 1358 -524
rect 1490 452 1536 464
rect 1490 -524 1496 452
rect 1530 -524 1536 452
rect 1490 -536 1536 -524
rect 1668 452 1714 464
rect 1668 -524 1674 452
rect 1708 -524 1714 452
rect 1668 -536 1714 -524
rect 1846 452 1892 464
rect 1846 -524 1852 452
rect 1886 -524 1892 452
rect 1846 -536 1892 -524
rect 2024 452 2070 464
rect 2024 -524 2030 452
rect 2064 -524 2070 452
rect 2024 -536 2070 -524
rect 2202 452 2248 464
rect 2202 -524 2208 452
rect 2242 -524 2248 452
rect 2202 -536 2248 -524
rect 2380 452 2426 464
rect 2380 -524 2386 452
rect 2420 -524 2426 452
rect 2380 -536 2426 -524
rect 2558 452 2604 464
rect 2558 -524 2564 452
rect 2598 -524 2604 452
rect 2558 -536 2604 -524
rect 2736 452 2782 464
rect 2736 -524 2742 452
rect 2776 -524 2782 452
rect 2736 -536 2782 -524
rect 2914 452 2960 464
rect 2914 -524 2920 452
rect 2954 -524 2960 452
rect 2914 -536 2960 -524
rect 3092 452 3138 464
rect 3092 -524 3098 452
rect 3132 -524 3138 452
rect 3092 -536 3138 -524
rect 3270 452 3316 464
rect 3270 -524 3276 452
rect 3310 -524 3316 452
rect 3270 -536 3316 -524
rect 3448 452 3494 464
rect 3448 -524 3454 452
rect 3488 -524 3494 452
rect 3448 -536 3494 -524
rect 3626 452 3672 464
rect 3626 -524 3632 452
rect 3666 -524 3672 452
rect 3626 -536 3672 -524
rect 3804 452 3850 464
rect 3804 -524 3810 452
rect 3844 -524 3850 452
rect 3804 -536 3850 -524
rect 3982 452 4028 464
rect 3982 -524 3988 452
rect 4022 -524 4028 452
rect 3982 -536 4028 -524
rect 4160 452 4206 464
rect 4160 -524 4166 452
rect 4200 -524 4206 452
rect 4160 -536 4206 -524
<< properties >>
string FIXED_BBOX -4317 -667 4317 667
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 47 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

* NGSPICE file created from brownout_dig.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

.subckt brownout_dig VGND VPWR brout_filt ena force_rc_osc force_short_oneshot osc_ck
+ osc_ena otrip[0] otrip[1] otrip[2] otrip_decoded[0] otrip_decoded[1] otrip_decoded[2]
+ otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6] otrip_decoded[7]
+ out_unbuf timed_out vtrip[0] vtrip[1] vtrip[2] vtrip_decoded[0] vtrip_decoded[1]
+ vtrip_decoded[2] vtrip_decoded[3] vtrip_decoded[4] vtrip_decoded[5] vtrip_decoded[6]
+ vtrip_decoded[7]
X_062_ net10 net9 net8 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__and3b_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_114_ clknet_1_1__leaf_osc_ck _010_ net33 VGND VGND VPWR VPWR cnt\[10\] sky130_fd_sc_hd__dfstp_1
X_045_ cnt\[1\] cnt\[0\] cnt\[3\] cnt\[2\] VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and4_1
Xoutput20 net20 VGND VGND VPWR VPWR out_unbuf sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_061_ net10 net8 net9 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nor3b_1
X_113_ clknet_1_1__leaf_osc_ck _009_ net33 VGND VGND VPWR VPWR cnt\[9\] sky130_fd_sc_hd__dfstp_1
X_044_ cnt\[1\] cnt\[0\] cnt\[2\] VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and3_1
X_116__32 VGND VGND VPWR VPWR net32 _116__32/LO sky130_fd_sc_hd__conb_1
Xoutput21 net21 VGND VGND VPWR VPWR timed_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_060_ net10 net9 net8 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_8_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_112_ clknet_1_1__leaf_osc_ck _008_ net31 VGND VGND VPWR VPWR cnt\[8\] sky130_fd_sc_hd__dfstp_1
X_043_ net2 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput11 net11 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput22 net22 VGND VGND VPWR VPWR vtrip_decoded[0] sky130_fd_sc_hd__buf_2
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_111_ clknet_1_1__leaf_osc_ck _007_ net31 VGND VGND VPWR VPWR cnt\[7\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_12_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ brout_filt_retimed VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput23 net23 VGND VGND VPWR VPWR vtrip_decoded[1] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ clknet_1_1__leaf_osc_ck _006_ net31 VGND VGND VPWR VPWR cnt\[6\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_15_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR vtrip_decoded[2] sky130_fd_sc_hd__buf_2
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput25 net25 VGND VGND VPWR VPWR vtrip_decoded[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
X_099_ _030_ net30 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__nand2_1
Xoutput26 net26 VGND VGND VPWR VPWR vtrip_decoded[4] sky130_fd_sc_hd__clkbuf_4
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ cnt\[9\] _029_ net30 cnt\[10\] VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput27 net27 VGND VGND VPWR VPWR vtrip_decoded[5] sky130_fd_sc_hd__clkbuf_4
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
XFILLER_0_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_097_ _024_ _018_ _019_ _031_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput28 net28 VGND VGND VPWR VPWR vtrip_decoded[6] sky130_fd_sc_hd__clkbuf_4
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout30 _041_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ cnt\[9\] _029_ net30 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_6_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR vtrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
X_079_ _033_ _037_ net36 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_095_ _029_ _041_ cnt\[9\] VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21o_1
Xfanout31 net33 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ cnt\[3\] _026_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_094_ _024_ _016_ _017_ _031_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_077_ _033_ _036_ net36 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_14_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ _029_ net30 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_076_ _026_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__or2_1
Xinput1 brout_filt VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_059_ net10 net9 net8 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ cnt\[7\] cnt\[6\] net30 cnt\[8\] VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a31o_1
Xinput2 ena VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_075_ cnt\[1\] cnt\[0\] cnt\[2\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ net7 net5 net6 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and3_1
X_091_ _024_ _014_ _015_ _031_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 force_rc_osc VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_074_ _033_ _034_ net36 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a21oi_1
X_057_ net5 net6 net7 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_109_ clknet_1_0__leaf_osc_ck _005_ net31 VGND VGND VPWR VPWR cnt\[5\] sky130_fd_sc_hd__dfstp_1
X_090_ cnt\[7\] cnt\[6\] net30 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_9_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 force_short_oneshot VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_056_ net6 net5 net7 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3b_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_073_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_3_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_108_ clknet_1_0__leaf_osc_ck _004_ net31 VGND VGND VPWR VPWR cnt\[4\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_072_ cnt\[0\] _033_ net36 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__a21oi_1
Xinput5 otrip[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_055_ net5 net6 net7 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__nor3b_1
X_107_ clknet_1_0__leaf_osc_ck _003_ net31 VGND VGND VPWR VPWR cnt\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_071_ cnt\[11\] _028_ _030_ net4 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a31oi_4
Xinput6 otrip[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
X_054_ net7 net5 net6 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_106_ clknet_1_0__leaf_osc_ck _002_ net31 VGND VGND VPWR VPWR cnt\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 otrip[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_070_ _025_ _031_ _032_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__o21ai_1
Xinput10 vtrip[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
X_053_ net7 net5 net6 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_4_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_105_ clknet_1_0__leaf_osc_ck _001_ net31 VGND VGND VPWR VPWR cnt\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
Xinput8 vtrip[0] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_11_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_104_ clknet_1_0__leaf_osc_ck _000_ net31 VGND VGND VPWR VPWR cnt\[0\] sky130_fd_sc_hd__dfstp_1
X_052_ net7 net6 net5 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor3b_1
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 vtrip[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_051_ net7 net5 net6 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor3_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_103_ _024_ _022_ _023_ _031_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 cnt_rsb VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_050_ _024_ net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and2_1
X_102_ cnt\[11\] _030_ _041_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__nand3_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
Xhold2 cnt_rsb_stg2 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ _030_ net30 cnt\[11\] VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a21o_1
Xhold3 cnt_rsb_stg1 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _024_ _020_ _021_ _031_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_7_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 brout_filt_retimed VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_5_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ cnt\[6\] net30 cnt\[7\] VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ _024_ _012_ _013_ _031_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_9_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ cnt\[6\] net30 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_086_ cnt\[6\] net30 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ net3 brout_filt_ena_rsb VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ cnt\[5\] cnt\[4\] _027_ net4 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_068_ net1 net2 VGND VGND VPWR VPWR brout_filt_ena_rsb sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_13_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_067_ _024_ cnt\[11\] _028_ _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and4_2
X_084_ _033_ _040_ net36 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_119_ clknet_1_0__leaf_osc_ck net1 brout_filt_ena_rsb VGND VGND VPWR VPWR brout_filt_retimed
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ _028_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_066_ net10 net9 net8 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__and3_1
X_049_ cnt\[11\] _028_ _030_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and3_1
X_118_ clknet_1_1__leaf_osc_ck net34 net2 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 otrip[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_065_ net8 net9 net10 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_12_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_082_ cnt\[4\] _027_ cnt\[5\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_048_ cnt\[9\] cnt\[10\] _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__and3_2
X_117_ clknet_1_0__leaf_osc_ck net35 net2 VGND VGND VPWR VPWR cnt_rsb_stg2 sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 otrip[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_081_ _033_ _038_ net36 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_064_ net9 net8 net10 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__and3b_1
XFILLER_0_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 vtrip[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ cnt\[7\] cnt\[6\] cnt\[8\] VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and3_1
X_116_ clknet_1_1__leaf_osc_ck net32 net2 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ net9 net8 net10 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__nor3b_1
X_080_ cnt\[4\] _027_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ clknet_1_1__leaf_osc_ck _011_ net31 VGND VGND VPWR VPWR cnt\[11\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_8_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_046_ cnt\[5\] cnt\[4\] _027_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and3_1
XANTENNA_4 vtrip[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends


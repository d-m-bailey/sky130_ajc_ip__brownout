magic
tech sky130A
magscale 1 2
timestamp 1712947988
<< pwell >>
rect -1463 -358 1463 358
<< mvnmos >>
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
<< mvndiff >>
rect -1293 88 -1235 100
rect -1293 -88 -1281 88
rect -1247 -88 -1235 88
rect -1293 -100 -1235 -88
rect -1135 88 -1077 100
rect -1135 -88 -1123 88
rect -1089 -88 -1077 88
rect -1135 -100 -1077 -88
rect -977 88 -919 100
rect -977 -88 -965 88
rect -931 -88 -919 88
rect -977 -100 -919 -88
rect -819 88 -761 100
rect -819 -88 -807 88
rect -773 -88 -761 88
rect -819 -100 -761 -88
rect -661 88 -603 100
rect -661 -88 -649 88
rect -615 -88 -603 88
rect -661 -100 -603 -88
rect -503 88 -445 100
rect -503 -88 -491 88
rect -457 -88 -445 88
rect -503 -100 -445 -88
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
rect 445 88 503 100
rect 445 -88 457 88
rect 491 -88 503 88
rect 445 -100 503 -88
rect 603 88 661 100
rect 603 -88 615 88
rect 649 -88 661 88
rect 603 -100 661 -88
rect 761 88 819 100
rect 761 -88 773 88
rect 807 -88 819 88
rect 761 -100 819 -88
rect 919 88 977 100
rect 919 -88 931 88
rect 965 -88 977 88
rect 919 -100 977 -88
rect 1077 88 1135 100
rect 1077 -88 1089 88
rect 1123 -88 1135 88
rect 1077 -100 1135 -88
rect 1235 88 1293 100
rect 1235 -88 1247 88
rect 1281 -88 1293 88
rect 1235 -100 1293 -88
<< mvndiffc >>
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
<< mvpsubdiff >>
rect -1427 310 1427 322
rect -1427 276 -1319 310
rect 1319 276 1427 310
rect -1427 264 1427 276
rect -1427 214 -1369 264
rect -1427 -214 -1415 214
rect -1381 -214 -1369 214
rect 1369 214 1427 264
rect -1427 -264 -1369 -214
rect 1369 -214 1381 214
rect 1415 -214 1427 214
rect 1369 -264 1427 -214
rect -1427 -276 1427 -264
rect -1427 -310 -1319 -276
rect 1319 -310 1427 -276
rect -1427 -322 1427 -310
<< mvpsubdiffcont >>
rect -1319 276 1319 310
rect -1415 -214 -1381 214
rect 1381 -214 1415 214
rect -1319 -310 1319 -276
<< poly >>
rect -1235 172 -1135 188
rect -1235 138 -1219 172
rect -1151 138 -1135 172
rect -1235 100 -1135 138
rect -1077 172 -977 188
rect -1077 138 -1061 172
rect -993 138 -977 172
rect -1077 100 -977 138
rect -919 172 -819 188
rect -919 138 -903 172
rect -835 138 -819 172
rect -919 100 -819 138
rect -761 172 -661 188
rect -761 138 -745 172
rect -677 138 -661 172
rect -761 100 -661 138
rect -603 172 -503 188
rect -603 138 -587 172
rect -519 138 -503 172
rect -603 100 -503 138
rect -445 172 -345 188
rect -445 138 -429 172
rect -361 138 -345 172
rect -445 100 -345 138
rect -287 172 -187 188
rect -287 138 -271 172
rect -203 138 -187 172
rect -287 100 -187 138
rect -129 172 -29 188
rect -129 138 -113 172
rect -45 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 45 172
rect 113 138 129 172
rect 29 100 129 138
rect 187 172 287 188
rect 187 138 203 172
rect 271 138 287 172
rect 187 100 287 138
rect 345 172 445 188
rect 345 138 361 172
rect 429 138 445 172
rect 345 100 445 138
rect 503 172 603 188
rect 503 138 519 172
rect 587 138 603 172
rect 503 100 603 138
rect 661 172 761 188
rect 661 138 677 172
rect 745 138 761 172
rect 661 100 761 138
rect 819 172 919 188
rect 819 138 835 172
rect 903 138 919 172
rect 819 100 919 138
rect 977 172 1077 188
rect 977 138 993 172
rect 1061 138 1077 172
rect 977 100 1077 138
rect 1135 172 1235 188
rect 1135 138 1151 172
rect 1219 138 1235 172
rect 1135 100 1235 138
rect -1235 -138 -1135 -100
rect -1235 -172 -1219 -138
rect -1151 -172 -1135 -138
rect -1235 -188 -1135 -172
rect -1077 -138 -977 -100
rect -1077 -172 -1061 -138
rect -993 -172 -977 -138
rect -1077 -188 -977 -172
rect -919 -138 -819 -100
rect -919 -172 -903 -138
rect -835 -172 -819 -138
rect -919 -188 -819 -172
rect -761 -138 -661 -100
rect -761 -172 -745 -138
rect -677 -172 -661 -138
rect -761 -188 -661 -172
rect -603 -138 -503 -100
rect -603 -172 -587 -138
rect -519 -172 -503 -138
rect -603 -188 -503 -172
rect -445 -138 -345 -100
rect -445 -172 -429 -138
rect -361 -172 -345 -138
rect -445 -188 -345 -172
rect -287 -138 -187 -100
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -287 -188 -187 -172
rect -129 -138 -29 -100
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 29 -188 129 -172
rect 187 -138 287 -100
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 187 -188 287 -172
rect 345 -138 445 -100
rect 345 -172 361 -138
rect 429 -172 445 -138
rect 345 -188 445 -172
rect 503 -138 603 -100
rect 503 -172 519 -138
rect 587 -172 603 -138
rect 503 -188 603 -172
rect 661 -138 761 -100
rect 661 -172 677 -138
rect 745 -172 761 -138
rect 661 -188 761 -172
rect 819 -138 919 -100
rect 819 -172 835 -138
rect 903 -172 919 -138
rect 819 -188 919 -172
rect 977 -138 1077 -100
rect 977 -172 993 -138
rect 1061 -172 1077 -138
rect 977 -188 1077 -172
rect 1135 -138 1235 -100
rect 1135 -172 1151 -138
rect 1219 -172 1235 -138
rect 1135 -188 1235 -172
<< polycont >>
rect -1219 138 -1151 172
rect -1061 138 -993 172
rect -903 138 -835 172
rect -745 138 -677 172
rect -587 138 -519 172
rect -429 138 -361 172
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect 361 138 429 172
rect 519 138 587 172
rect 677 138 745 172
rect 835 138 903 172
rect 993 138 1061 172
rect 1151 138 1219 172
rect -1219 -172 -1151 -138
rect -1061 -172 -993 -138
rect -903 -172 -835 -138
rect -745 -172 -677 -138
rect -587 -172 -519 -138
rect -429 -172 -361 -138
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
rect 361 -172 429 -138
rect 519 -172 587 -138
rect 677 -172 745 -138
rect 835 -172 903 -138
rect 993 -172 1061 -138
rect 1151 -172 1219 -138
<< locali >>
rect -1415 276 -1319 310
rect 1319 276 1415 310
rect -1415 214 -1381 276
rect 1381 214 1415 276
rect -1235 138 -1219 172
rect -1151 138 -1135 172
rect -1077 138 -1061 172
rect -993 138 -977 172
rect -919 138 -903 172
rect -835 138 -819 172
rect -761 138 -745 172
rect -677 138 -661 172
rect -603 138 -587 172
rect -519 138 -503 172
rect -445 138 -429 172
rect -361 138 -345 172
rect -287 138 -271 172
rect -203 138 -187 172
rect -129 138 -113 172
rect -45 138 -29 172
rect 29 138 45 172
rect 113 138 129 172
rect 187 138 203 172
rect 271 138 287 172
rect 345 138 361 172
rect 429 138 445 172
rect 503 138 519 172
rect 587 138 603 172
rect 661 138 677 172
rect 745 138 761 172
rect 819 138 835 172
rect 903 138 919 172
rect 977 138 993 172
rect 1061 138 1077 172
rect 1135 138 1151 172
rect 1219 138 1235 172
rect -1281 88 -1247 104
rect -1281 -104 -1247 -88
rect -1123 88 -1089 104
rect -1123 -104 -1089 -88
rect -965 88 -931 104
rect -965 -104 -931 -88
rect -807 88 -773 104
rect -807 -104 -773 -88
rect -649 88 -615 104
rect -649 -104 -615 -88
rect -491 88 -457 104
rect -491 -104 -457 -88
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect 457 88 491 104
rect 457 -104 491 -88
rect 615 88 649 104
rect 615 -104 649 -88
rect 773 88 807 104
rect 773 -104 807 -88
rect 931 88 965 104
rect 931 -104 965 -88
rect 1089 88 1123 104
rect 1089 -104 1123 -88
rect 1247 88 1281 104
rect 1247 -104 1281 -88
rect -1235 -172 -1219 -138
rect -1151 -172 -1135 -138
rect -1077 -172 -1061 -138
rect -993 -172 -977 -138
rect -919 -172 -903 -138
rect -835 -172 -819 -138
rect -761 -172 -745 -138
rect -677 -172 -661 -138
rect -603 -172 -587 -138
rect -519 -172 -503 -138
rect -445 -172 -429 -138
rect -361 -172 -345 -138
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 345 -172 361 -138
rect 429 -172 445 -138
rect 503 -172 519 -138
rect 587 -172 603 -138
rect 661 -172 677 -138
rect 745 -172 761 -138
rect 819 -172 835 -138
rect 903 -172 919 -138
rect 977 -172 993 -138
rect 1061 -172 1077 -138
rect 1135 -172 1151 -138
rect 1219 -172 1235 -138
rect -1415 -276 -1381 -214
rect 1381 -276 1415 -214
rect -1415 -310 -1319 -276
rect 1319 -310 1415 -276
<< viali >>
rect -1219 138 -1151 172
rect -1061 138 -993 172
rect -903 138 -835 172
rect -745 138 -677 172
rect -587 138 -519 172
rect -429 138 -361 172
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect 361 138 429 172
rect 519 138 587 172
rect 677 138 745 172
rect 835 138 903 172
rect 993 138 1061 172
rect 1151 138 1219 172
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect -1219 -172 -1151 -138
rect -1061 -172 -993 -138
rect -903 -172 -835 -138
rect -745 -172 -677 -138
rect -587 -172 -519 -138
rect -429 -172 -361 -138
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
rect 361 -172 429 -138
rect 519 -172 587 -138
rect 677 -172 745 -138
rect 835 -172 903 -138
rect 993 -172 1061 -138
rect 1151 -172 1219 -138
<< metal1 >>
rect -1231 172 -1139 178
rect -1231 138 -1219 172
rect -1151 138 -1139 172
rect -1231 132 -1139 138
rect -1073 172 -981 178
rect -1073 138 -1061 172
rect -993 138 -981 172
rect -1073 132 -981 138
rect -915 172 -823 178
rect -915 138 -903 172
rect -835 138 -823 172
rect -915 132 -823 138
rect -757 172 -665 178
rect -757 138 -745 172
rect -677 138 -665 172
rect -757 132 -665 138
rect -599 172 -507 178
rect -599 138 -587 172
rect -519 138 -507 172
rect -599 132 -507 138
rect -441 172 -349 178
rect -441 138 -429 172
rect -361 138 -349 172
rect -441 132 -349 138
rect -283 172 -191 178
rect -283 138 -271 172
rect -203 138 -191 172
rect -283 132 -191 138
rect -125 172 -33 178
rect -125 138 -113 172
rect -45 138 -33 172
rect -125 132 -33 138
rect 33 172 125 178
rect 33 138 45 172
rect 113 138 125 172
rect 33 132 125 138
rect 191 172 283 178
rect 191 138 203 172
rect 271 138 283 172
rect 191 132 283 138
rect 349 172 441 178
rect 349 138 361 172
rect 429 138 441 172
rect 349 132 441 138
rect 507 172 599 178
rect 507 138 519 172
rect 587 138 599 172
rect 507 132 599 138
rect 665 172 757 178
rect 665 138 677 172
rect 745 138 757 172
rect 665 132 757 138
rect 823 172 915 178
rect 823 138 835 172
rect 903 138 915 172
rect 823 132 915 138
rect 981 172 1073 178
rect 981 138 993 172
rect 1061 138 1073 172
rect 981 132 1073 138
rect 1139 172 1231 178
rect 1139 138 1151 172
rect 1219 138 1231 172
rect 1139 132 1231 138
rect -1287 88 -1241 100
rect -1287 -88 -1281 88
rect -1247 -88 -1241 88
rect -1287 -100 -1241 -88
rect -1129 88 -1083 100
rect -1129 -88 -1123 88
rect -1089 -88 -1083 88
rect -1129 -100 -1083 -88
rect -971 88 -925 100
rect -971 -88 -965 88
rect -931 -88 -925 88
rect -971 -100 -925 -88
rect -813 88 -767 100
rect -813 -88 -807 88
rect -773 -88 -767 88
rect -813 -100 -767 -88
rect -655 88 -609 100
rect -655 -88 -649 88
rect -615 -88 -609 88
rect -655 -100 -609 -88
rect -497 88 -451 100
rect -497 -88 -491 88
rect -457 -88 -451 88
rect -497 -100 -451 -88
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect 451 88 497 100
rect 451 -88 457 88
rect 491 -88 497 88
rect 451 -100 497 -88
rect 609 88 655 100
rect 609 -88 615 88
rect 649 -88 655 88
rect 609 -100 655 -88
rect 767 88 813 100
rect 767 -88 773 88
rect 807 -88 813 88
rect 767 -100 813 -88
rect 925 88 971 100
rect 925 -88 931 88
rect 965 -88 971 88
rect 925 -100 971 -88
rect 1083 88 1129 100
rect 1083 -88 1089 88
rect 1123 -88 1129 88
rect 1083 -100 1129 -88
rect 1241 88 1287 100
rect 1241 -88 1247 88
rect 1281 -88 1287 88
rect 1241 -100 1287 -88
rect -1231 -138 -1139 -132
rect -1231 -172 -1219 -138
rect -1151 -172 -1139 -138
rect -1231 -178 -1139 -172
rect -1073 -138 -981 -132
rect -1073 -172 -1061 -138
rect -993 -172 -981 -138
rect -1073 -178 -981 -172
rect -915 -138 -823 -132
rect -915 -172 -903 -138
rect -835 -172 -823 -138
rect -915 -178 -823 -172
rect -757 -138 -665 -132
rect -757 -172 -745 -138
rect -677 -172 -665 -138
rect -757 -178 -665 -172
rect -599 -138 -507 -132
rect -599 -172 -587 -138
rect -519 -172 -507 -138
rect -599 -178 -507 -172
rect -441 -138 -349 -132
rect -441 -172 -429 -138
rect -361 -172 -349 -138
rect -441 -178 -349 -172
rect -283 -138 -191 -132
rect -283 -172 -271 -138
rect -203 -172 -191 -138
rect -283 -178 -191 -172
rect -125 -138 -33 -132
rect -125 -172 -113 -138
rect -45 -172 -33 -138
rect -125 -178 -33 -172
rect 33 -138 125 -132
rect 33 -172 45 -138
rect 113 -172 125 -138
rect 33 -178 125 -172
rect 191 -138 283 -132
rect 191 -172 203 -138
rect 271 -172 283 -138
rect 191 -178 283 -172
rect 349 -138 441 -132
rect 349 -172 361 -138
rect 429 -172 441 -138
rect 349 -178 441 -172
rect 507 -138 599 -132
rect 507 -172 519 -138
rect 587 -172 599 -138
rect 507 -178 599 -172
rect 665 -138 757 -132
rect 665 -172 677 -138
rect 745 -172 757 -138
rect 665 -178 757 -172
rect 823 -138 915 -132
rect 823 -172 835 -138
rect 903 -172 915 -138
rect 823 -178 915 -172
rect 981 -138 1073 -132
rect 981 -172 993 -138
rect 1061 -172 1073 -138
rect 981 -178 1073 -172
rect 1139 -138 1231 -132
rect 1139 -172 1151 -138
rect 1219 -172 1231 -138
rect 1139 -178 1231 -172
<< properties >>
string FIXED_BBOX -1398 -293 1398 293
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

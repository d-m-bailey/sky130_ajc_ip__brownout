magic
tech sky130A
magscale 1 2
timestamp 1712930986
<< pwell >>
rect -328 -1039 328 1039
<< mvnmos >>
rect -100 581 100 781
rect -100 225 100 425
rect -100 -131 100 69
rect -100 -487 100 -287
rect -100 -843 100 -643
<< mvndiff >>
rect -158 769 -100 781
rect -158 593 -146 769
rect -112 593 -100 769
rect -158 581 -100 593
rect 100 769 158 781
rect 100 593 112 769
rect 146 593 158 769
rect 100 581 158 593
rect -158 413 -100 425
rect -158 237 -146 413
rect -112 237 -100 413
rect -158 225 -100 237
rect 100 413 158 425
rect 100 237 112 413
rect 146 237 158 413
rect 100 225 158 237
rect -158 57 -100 69
rect -158 -119 -146 57
rect -112 -119 -100 57
rect -158 -131 -100 -119
rect 100 57 158 69
rect 100 -119 112 57
rect 146 -119 158 57
rect 100 -131 158 -119
rect -158 -299 -100 -287
rect -158 -475 -146 -299
rect -112 -475 -100 -299
rect -158 -487 -100 -475
rect 100 -299 158 -287
rect 100 -475 112 -299
rect 146 -475 158 -299
rect 100 -487 158 -475
rect -158 -655 -100 -643
rect -158 -831 -146 -655
rect -112 -831 -100 -655
rect -158 -843 -100 -831
rect 100 -655 158 -643
rect 100 -831 112 -655
rect 146 -831 158 -655
rect 100 -843 158 -831
<< mvndiffc >>
rect -146 593 -112 769
rect 112 593 146 769
rect -146 237 -112 413
rect 112 237 146 413
rect -146 -119 -112 57
rect 112 -119 146 57
rect -146 -475 -112 -299
rect 112 -475 146 -299
rect -146 -831 -112 -655
rect 112 -831 146 -655
<< mvpsubdiff >>
rect -292 991 292 1003
rect -292 957 -184 991
rect 184 957 292 991
rect -292 945 292 957
rect -292 895 -234 945
rect -292 -895 -280 895
rect -246 -895 -234 895
rect 234 895 292 945
rect -292 -945 -234 -895
rect 234 -895 246 895
rect 280 -895 292 895
rect 234 -945 292 -895
rect -292 -957 292 -945
rect -292 -991 -184 -957
rect 184 -991 292 -957
rect -292 -1003 292 -991
<< mvpsubdiffcont >>
rect -184 957 184 991
rect -280 -895 -246 895
rect 246 -895 280 895
rect -184 -991 184 -957
<< poly >>
rect -100 853 100 869
rect -100 819 -84 853
rect 84 819 100 853
rect -100 781 100 819
rect -100 555 100 581
rect -100 497 100 513
rect -100 463 -84 497
rect 84 463 100 497
rect -100 425 100 463
rect -100 199 100 225
rect -100 141 100 157
rect -100 107 -84 141
rect 84 107 100 141
rect -100 69 100 107
rect -100 -157 100 -131
rect -100 -215 100 -199
rect -100 -249 -84 -215
rect 84 -249 100 -215
rect -100 -287 100 -249
rect -100 -513 100 -487
rect -100 -571 100 -555
rect -100 -605 -84 -571
rect 84 -605 100 -571
rect -100 -643 100 -605
rect -100 -869 100 -843
<< polycont >>
rect -84 819 84 853
rect -84 463 84 497
rect -84 107 84 141
rect -84 -249 84 -215
rect -84 -605 84 -571
<< locali >>
rect -280 957 -184 991
rect 184 957 280 991
rect -280 895 -246 957
rect 246 895 280 957
rect -100 819 -84 853
rect 84 819 100 853
rect -146 769 -112 785
rect -146 577 -112 593
rect 112 769 146 785
rect 112 577 146 593
rect -100 463 -84 497
rect 84 463 100 497
rect -146 413 -112 429
rect -146 221 -112 237
rect 112 413 146 429
rect 112 221 146 237
rect -100 107 -84 141
rect 84 107 100 141
rect -146 57 -112 73
rect -146 -135 -112 -119
rect 112 57 146 73
rect 112 -135 146 -119
rect -100 -249 -84 -215
rect 84 -249 100 -215
rect -146 -299 -112 -283
rect -146 -491 -112 -475
rect 112 -299 146 -283
rect 112 -491 146 -475
rect -100 -605 -84 -571
rect 84 -605 100 -571
rect -146 -655 -112 -639
rect -146 -847 -112 -831
rect 112 -655 146 -639
rect 112 -847 146 -831
rect -280 -957 -246 -895
rect 246 -957 280 -895
rect -280 -991 -184 -957
rect 184 -991 280 -957
<< viali >>
rect -84 819 84 853
rect -146 593 -112 769
rect 112 593 146 769
rect -84 463 84 497
rect -146 237 -112 413
rect 112 237 146 413
rect -84 107 84 141
rect -146 -119 -112 57
rect 112 -119 146 57
rect -84 -249 84 -215
rect -146 -475 -112 -299
rect 112 -475 146 -299
rect -84 -605 84 -571
rect -146 -831 -112 -655
rect 112 -831 146 -655
<< metal1 >>
rect -96 853 96 859
rect -96 819 -84 853
rect 84 819 96 853
rect -96 813 96 819
rect -152 769 -106 781
rect -152 593 -146 769
rect -112 593 -106 769
rect -152 581 -106 593
rect 106 769 152 781
rect 106 593 112 769
rect 146 593 152 769
rect 106 581 152 593
rect -96 497 96 503
rect -96 463 -84 497
rect 84 463 96 497
rect -96 457 96 463
rect -152 413 -106 425
rect -152 237 -146 413
rect -112 237 -106 413
rect -152 225 -106 237
rect 106 413 152 425
rect 106 237 112 413
rect 146 237 152 413
rect 106 225 152 237
rect -96 141 96 147
rect -96 107 -84 141
rect 84 107 96 141
rect -96 101 96 107
rect -152 57 -106 69
rect -152 -119 -146 57
rect -112 -119 -106 57
rect -152 -131 -106 -119
rect 106 57 152 69
rect 106 -119 112 57
rect 146 -119 152 57
rect 106 -131 152 -119
rect -96 -215 96 -209
rect -96 -249 -84 -215
rect 84 -249 96 -215
rect -96 -255 96 -249
rect -152 -299 -106 -287
rect -152 -475 -146 -299
rect -112 -475 -106 -299
rect -152 -487 -106 -475
rect 106 -299 152 -287
rect 106 -475 112 -299
rect 146 -475 152 -299
rect 106 -487 152 -475
rect -96 -571 96 -565
rect -96 -605 -84 -571
rect 84 -605 96 -571
rect -96 -611 96 -605
rect -152 -655 -106 -643
rect -152 -831 -146 -655
rect -112 -831 -106 -655
rect -152 -843 -106 -831
rect 106 -655 152 -643
rect 106 -831 112 -655
rect 146 -831 152 -655
rect 106 -843 152 -831
<< properties >>
string FIXED_BBOX -263 -974 263 974
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

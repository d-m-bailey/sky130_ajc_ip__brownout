magic
tech sky130A
magscale 1 2
timestamp 1712722749
<< nwell >>
rect -452 -164 452 198
<< pmos >>
rect -358 -64 -158 136
rect -100 -64 100 136
rect 158 -64 358 136
<< pdiff >>
rect -416 124 -358 136
rect -416 -52 -404 124
rect -370 -52 -358 124
rect -416 -64 -358 -52
rect -158 124 -100 136
rect -158 -52 -146 124
rect -112 -52 -100 124
rect -158 -64 -100 -52
rect 100 124 158 136
rect 100 -52 112 124
rect 146 -52 158 124
rect 100 -64 158 -52
rect 358 124 416 136
rect 358 -52 370 124
rect 404 -52 416 124
rect 358 -64 416 -52
<< pdiffc >>
rect -404 -52 -370 124
rect -146 -52 -112 124
rect 112 -52 146 124
rect 370 -52 404 124
<< poly >>
rect -358 136 -158 162
rect -100 136 100 162
rect 158 136 358 162
rect -358 -111 -158 -64
rect -358 -145 -342 -111
rect -174 -145 -158 -111
rect -358 -161 -158 -145
rect -100 -111 100 -64
rect -100 -145 -84 -111
rect 84 -145 100 -111
rect -100 -161 100 -145
rect 158 -111 358 -64
rect 158 -145 174 -111
rect 342 -145 358 -111
rect 158 -161 358 -145
<< polycont >>
rect -342 -145 -174 -111
rect -84 -145 84 -111
rect 174 -145 342 -111
<< locali >>
rect -404 124 -370 140
rect -404 -68 -370 -52
rect -146 124 -112 140
rect -146 -68 -112 -52
rect 112 124 146 140
rect 112 -68 146 -52
rect 370 124 404 140
rect 370 -68 404 -52
rect -358 -145 -342 -111
rect -174 -145 -158 -111
rect -100 -145 -84 -111
rect 84 -145 100 -111
rect 158 -145 174 -111
rect 342 -145 358 -111
<< viali >>
rect -404 -52 -370 124
rect -146 -52 -112 124
rect 112 -52 146 124
rect 370 -52 404 124
rect -342 -145 -174 -111
rect -84 -145 84 -111
rect 174 -145 342 -111
<< metal1 >>
rect -410 124 -364 136
rect -410 -52 -404 124
rect -370 -52 -364 124
rect -410 -64 -364 -52
rect -152 124 -106 136
rect -152 -52 -146 124
rect -112 -52 -106 124
rect -152 -64 -106 -52
rect 106 124 152 136
rect 106 -52 112 124
rect 146 -52 152 124
rect 106 -64 152 -52
rect 364 124 410 136
rect 364 -52 370 124
rect 404 -52 410 124
rect 364 -64 410 -52
rect -354 -111 -162 -105
rect -354 -145 -342 -111
rect -174 -145 -162 -111
rect -354 -151 -162 -145
rect -96 -111 96 -105
rect -96 -145 -84 -111
rect 84 -145 96 -111
rect -96 -151 96 -145
rect 162 -111 354 -105
rect 162 -145 174 -111
rect 342 -145 354 -111
rect 162 -151 354 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712543064
<< pwell >>
rect -3483 -1773 3483 1773
<< nmos >>
rect -3287 1363 -1687 1563
rect -1629 1363 -29 1563
rect 29 1363 1629 1563
rect 1687 1363 3287 1563
rect -3287 945 -1687 1145
rect -1629 945 -29 1145
rect 29 945 1629 1145
rect 1687 945 3287 1145
rect -3287 527 -1687 727
rect -1629 527 -29 727
rect 29 527 1629 727
rect 1687 527 3287 727
rect -3287 109 -1687 309
rect -1629 109 -29 309
rect 29 109 1629 309
rect 1687 109 3287 309
rect -3287 -309 -1687 -109
rect -1629 -309 -29 -109
rect 29 -309 1629 -109
rect 1687 -309 3287 -109
rect -3287 -727 -1687 -527
rect -1629 -727 -29 -527
rect 29 -727 1629 -527
rect 1687 -727 3287 -527
rect -3287 -1145 -1687 -945
rect -1629 -1145 -29 -945
rect 29 -1145 1629 -945
rect 1687 -1145 3287 -945
rect -3287 -1563 -1687 -1363
rect -1629 -1563 -29 -1363
rect 29 -1563 1629 -1363
rect 1687 -1563 3287 -1363
<< ndiff >>
rect -3345 1551 -3287 1563
rect -3345 1375 -3333 1551
rect -3299 1375 -3287 1551
rect -3345 1363 -3287 1375
rect -1687 1551 -1629 1563
rect -1687 1375 -1675 1551
rect -1641 1375 -1629 1551
rect -1687 1363 -1629 1375
rect -29 1551 29 1563
rect -29 1375 -17 1551
rect 17 1375 29 1551
rect -29 1363 29 1375
rect 1629 1551 1687 1563
rect 1629 1375 1641 1551
rect 1675 1375 1687 1551
rect 1629 1363 1687 1375
rect 3287 1551 3345 1563
rect 3287 1375 3299 1551
rect 3333 1375 3345 1551
rect 3287 1363 3345 1375
rect -3345 1133 -3287 1145
rect -3345 957 -3333 1133
rect -3299 957 -3287 1133
rect -3345 945 -3287 957
rect -1687 1133 -1629 1145
rect -1687 957 -1675 1133
rect -1641 957 -1629 1133
rect -1687 945 -1629 957
rect -29 1133 29 1145
rect -29 957 -17 1133
rect 17 957 29 1133
rect -29 945 29 957
rect 1629 1133 1687 1145
rect 1629 957 1641 1133
rect 1675 957 1687 1133
rect 1629 945 1687 957
rect 3287 1133 3345 1145
rect 3287 957 3299 1133
rect 3333 957 3345 1133
rect 3287 945 3345 957
rect -3345 715 -3287 727
rect -3345 539 -3333 715
rect -3299 539 -3287 715
rect -3345 527 -3287 539
rect -1687 715 -1629 727
rect -1687 539 -1675 715
rect -1641 539 -1629 715
rect -1687 527 -1629 539
rect -29 715 29 727
rect -29 539 -17 715
rect 17 539 29 715
rect -29 527 29 539
rect 1629 715 1687 727
rect 1629 539 1641 715
rect 1675 539 1687 715
rect 1629 527 1687 539
rect 3287 715 3345 727
rect 3287 539 3299 715
rect 3333 539 3345 715
rect 3287 527 3345 539
rect -3345 297 -3287 309
rect -3345 121 -3333 297
rect -3299 121 -3287 297
rect -3345 109 -3287 121
rect -1687 297 -1629 309
rect -1687 121 -1675 297
rect -1641 121 -1629 297
rect -1687 109 -1629 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 1629 297 1687 309
rect 1629 121 1641 297
rect 1675 121 1687 297
rect 1629 109 1687 121
rect 3287 297 3345 309
rect 3287 121 3299 297
rect 3333 121 3345 297
rect 3287 109 3345 121
rect -3345 -121 -3287 -109
rect -3345 -297 -3333 -121
rect -3299 -297 -3287 -121
rect -3345 -309 -3287 -297
rect -1687 -121 -1629 -109
rect -1687 -297 -1675 -121
rect -1641 -297 -1629 -121
rect -1687 -309 -1629 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 1629 -121 1687 -109
rect 1629 -297 1641 -121
rect 1675 -297 1687 -121
rect 1629 -309 1687 -297
rect 3287 -121 3345 -109
rect 3287 -297 3299 -121
rect 3333 -297 3345 -121
rect 3287 -309 3345 -297
rect -3345 -539 -3287 -527
rect -3345 -715 -3333 -539
rect -3299 -715 -3287 -539
rect -3345 -727 -3287 -715
rect -1687 -539 -1629 -527
rect -1687 -715 -1675 -539
rect -1641 -715 -1629 -539
rect -1687 -727 -1629 -715
rect -29 -539 29 -527
rect -29 -715 -17 -539
rect 17 -715 29 -539
rect -29 -727 29 -715
rect 1629 -539 1687 -527
rect 1629 -715 1641 -539
rect 1675 -715 1687 -539
rect 1629 -727 1687 -715
rect 3287 -539 3345 -527
rect 3287 -715 3299 -539
rect 3333 -715 3345 -539
rect 3287 -727 3345 -715
rect -3345 -957 -3287 -945
rect -3345 -1133 -3333 -957
rect -3299 -1133 -3287 -957
rect -3345 -1145 -3287 -1133
rect -1687 -957 -1629 -945
rect -1687 -1133 -1675 -957
rect -1641 -1133 -1629 -957
rect -1687 -1145 -1629 -1133
rect -29 -957 29 -945
rect -29 -1133 -17 -957
rect 17 -1133 29 -957
rect -29 -1145 29 -1133
rect 1629 -957 1687 -945
rect 1629 -1133 1641 -957
rect 1675 -1133 1687 -957
rect 1629 -1145 1687 -1133
rect 3287 -957 3345 -945
rect 3287 -1133 3299 -957
rect 3333 -1133 3345 -957
rect 3287 -1145 3345 -1133
rect -3345 -1375 -3287 -1363
rect -3345 -1551 -3333 -1375
rect -3299 -1551 -3287 -1375
rect -3345 -1563 -3287 -1551
rect -1687 -1375 -1629 -1363
rect -1687 -1551 -1675 -1375
rect -1641 -1551 -1629 -1375
rect -1687 -1563 -1629 -1551
rect -29 -1375 29 -1363
rect -29 -1551 -17 -1375
rect 17 -1551 29 -1375
rect -29 -1563 29 -1551
rect 1629 -1375 1687 -1363
rect 1629 -1551 1641 -1375
rect 1675 -1551 1687 -1375
rect 1629 -1563 1687 -1551
rect 3287 -1375 3345 -1363
rect 3287 -1551 3299 -1375
rect 3333 -1551 3345 -1375
rect 3287 -1563 3345 -1551
<< ndiffc >>
rect -3333 1375 -3299 1551
rect -1675 1375 -1641 1551
rect -17 1375 17 1551
rect 1641 1375 1675 1551
rect 3299 1375 3333 1551
rect -3333 957 -3299 1133
rect -1675 957 -1641 1133
rect -17 957 17 1133
rect 1641 957 1675 1133
rect 3299 957 3333 1133
rect -3333 539 -3299 715
rect -1675 539 -1641 715
rect -17 539 17 715
rect 1641 539 1675 715
rect 3299 539 3333 715
rect -3333 121 -3299 297
rect -1675 121 -1641 297
rect -17 121 17 297
rect 1641 121 1675 297
rect 3299 121 3333 297
rect -3333 -297 -3299 -121
rect -1675 -297 -1641 -121
rect -17 -297 17 -121
rect 1641 -297 1675 -121
rect 3299 -297 3333 -121
rect -3333 -715 -3299 -539
rect -1675 -715 -1641 -539
rect -17 -715 17 -539
rect 1641 -715 1675 -539
rect 3299 -715 3333 -539
rect -3333 -1133 -3299 -957
rect -1675 -1133 -1641 -957
rect -17 -1133 17 -957
rect 1641 -1133 1675 -957
rect 3299 -1133 3333 -957
rect -3333 -1551 -3299 -1375
rect -1675 -1551 -1641 -1375
rect -17 -1551 17 -1375
rect 1641 -1551 1675 -1375
rect 3299 -1551 3333 -1375
<< psubdiff >>
rect -3447 1703 -3351 1737
rect 3351 1703 3447 1737
rect -3447 1641 -3413 1703
rect 3413 1641 3447 1703
rect -3447 -1703 -3413 -1641
rect 3413 -1703 3447 -1641
rect -3447 -1737 -3351 -1703
rect 3351 -1737 3447 -1703
<< psubdiffcont >>
rect -3351 1703 3351 1737
rect -3447 -1641 -3413 1641
rect 3413 -1641 3447 1641
rect -3351 -1737 3351 -1703
<< poly >>
rect -3287 1635 -1687 1651
rect -3287 1601 -3271 1635
rect -1703 1601 -1687 1635
rect -3287 1563 -1687 1601
rect -1629 1635 -29 1651
rect -1629 1601 -1613 1635
rect -45 1601 -29 1635
rect -1629 1563 -29 1601
rect 29 1635 1629 1651
rect 29 1601 45 1635
rect 1613 1601 1629 1635
rect 29 1563 1629 1601
rect 1687 1635 3287 1651
rect 1687 1601 1703 1635
rect 3271 1601 3287 1635
rect 1687 1563 3287 1601
rect -3287 1325 -1687 1363
rect -3287 1291 -3271 1325
rect -1703 1291 -1687 1325
rect -3287 1275 -1687 1291
rect -1629 1325 -29 1363
rect -1629 1291 -1613 1325
rect -45 1291 -29 1325
rect -1629 1275 -29 1291
rect 29 1325 1629 1363
rect 29 1291 45 1325
rect 1613 1291 1629 1325
rect 29 1275 1629 1291
rect 1687 1325 3287 1363
rect 1687 1291 1703 1325
rect 3271 1291 3287 1325
rect 1687 1275 3287 1291
rect -3287 1217 -1687 1233
rect -3287 1183 -3271 1217
rect -1703 1183 -1687 1217
rect -3287 1145 -1687 1183
rect -1629 1217 -29 1233
rect -1629 1183 -1613 1217
rect -45 1183 -29 1217
rect -1629 1145 -29 1183
rect 29 1217 1629 1233
rect 29 1183 45 1217
rect 1613 1183 1629 1217
rect 29 1145 1629 1183
rect 1687 1217 3287 1233
rect 1687 1183 1703 1217
rect 3271 1183 3287 1217
rect 1687 1145 3287 1183
rect -3287 907 -1687 945
rect -3287 873 -3271 907
rect -1703 873 -1687 907
rect -3287 857 -1687 873
rect -1629 907 -29 945
rect -1629 873 -1613 907
rect -45 873 -29 907
rect -1629 857 -29 873
rect 29 907 1629 945
rect 29 873 45 907
rect 1613 873 1629 907
rect 29 857 1629 873
rect 1687 907 3287 945
rect 1687 873 1703 907
rect 3271 873 3287 907
rect 1687 857 3287 873
rect -3287 799 -1687 815
rect -3287 765 -3271 799
rect -1703 765 -1687 799
rect -3287 727 -1687 765
rect -1629 799 -29 815
rect -1629 765 -1613 799
rect -45 765 -29 799
rect -1629 727 -29 765
rect 29 799 1629 815
rect 29 765 45 799
rect 1613 765 1629 799
rect 29 727 1629 765
rect 1687 799 3287 815
rect 1687 765 1703 799
rect 3271 765 3287 799
rect 1687 727 3287 765
rect -3287 489 -1687 527
rect -3287 455 -3271 489
rect -1703 455 -1687 489
rect -3287 439 -1687 455
rect -1629 489 -29 527
rect -1629 455 -1613 489
rect -45 455 -29 489
rect -1629 439 -29 455
rect 29 489 1629 527
rect 29 455 45 489
rect 1613 455 1629 489
rect 29 439 1629 455
rect 1687 489 3287 527
rect 1687 455 1703 489
rect 3271 455 3287 489
rect 1687 439 3287 455
rect -3287 381 -1687 397
rect -3287 347 -3271 381
rect -1703 347 -1687 381
rect -3287 309 -1687 347
rect -1629 381 -29 397
rect -1629 347 -1613 381
rect -45 347 -29 381
rect -1629 309 -29 347
rect 29 381 1629 397
rect 29 347 45 381
rect 1613 347 1629 381
rect 29 309 1629 347
rect 1687 381 3287 397
rect 1687 347 1703 381
rect 3271 347 3287 381
rect 1687 309 3287 347
rect -3287 71 -1687 109
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -3287 21 -1687 37
rect -1629 71 -29 109
rect -1629 37 -1613 71
rect -45 37 -29 71
rect -1629 21 -29 37
rect 29 71 1629 109
rect 29 37 45 71
rect 1613 37 1629 71
rect 29 21 1629 37
rect 1687 71 3287 109
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 1687 21 3287 37
rect -3287 -37 -1687 -21
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -3287 -109 -1687 -71
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -109 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -109 1629 -71
rect 1687 -37 3287 -21
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 1687 -109 3287 -71
rect -3287 -347 -1687 -309
rect -3287 -381 -3271 -347
rect -1703 -381 -1687 -347
rect -3287 -397 -1687 -381
rect -1629 -347 -29 -309
rect -1629 -381 -1613 -347
rect -45 -381 -29 -347
rect -1629 -397 -29 -381
rect 29 -347 1629 -309
rect 29 -381 45 -347
rect 1613 -381 1629 -347
rect 29 -397 1629 -381
rect 1687 -347 3287 -309
rect 1687 -381 1703 -347
rect 3271 -381 3287 -347
rect 1687 -397 3287 -381
rect -3287 -455 -1687 -439
rect -3287 -489 -3271 -455
rect -1703 -489 -1687 -455
rect -3287 -527 -1687 -489
rect -1629 -455 -29 -439
rect -1629 -489 -1613 -455
rect -45 -489 -29 -455
rect -1629 -527 -29 -489
rect 29 -455 1629 -439
rect 29 -489 45 -455
rect 1613 -489 1629 -455
rect 29 -527 1629 -489
rect 1687 -455 3287 -439
rect 1687 -489 1703 -455
rect 3271 -489 3287 -455
rect 1687 -527 3287 -489
rect -3287 -765 -1687 -727
rect -3287 -799 -3271 -765
rect -1703 -799 -1687 -765
rect -3287 -815 -1687 -799
rect -1629 -765 -29 -727
rect -1629 -799 -1613 -765
rect -45 -799 -29 -765
rect -1629 -815 -29 -799
rect 29 -765 1629 -727
rect 29 -799 45 -765
rect 1613 -799 1629 -765
rect 29 -815 1629 -799
rect 1687 -765 3287 -727
rect 1687 -799 1703 -765
rect 3271 -799 3287 -765
rect 1687 -815 3287 -799
rect -3287 -873 -1687 -857
rect -3287 -907 -3271 -873
rect -1703 -907 -1687 -873
rect -3287 -945 -1687 -907
rect -1629 -873 -29 -857
rect -1629 -907 -1613 -873
rect -45 -907 -29 -873
rect -1629 -945 -29 -907
rect 29 -873 1629 -857
rect 29 -907 45 -873
rect 1613 -907 1629 -873
rect 29 -945 1629 -907
rect 1687 -873 3287 -857
rect 1687 -907 1703 -873
rect 3271 -907 3287 -873
rect 1687 -945 3287 -907
rect -3287 -1183 -1687 -1145
rect -3287 -1217 -3271 -1183
rect -1703 -1217 -1687 -1183
rect -3287 -1233 -1687 -1217
rect -1629 -1183 -29 -1145
rect -1629 -1217 -1613 -1183
rect -45 -1217 -29 -1183
rect -1629 -1233 -29 -1217
rect 29 -1183 1629 -1145
rect 29 -1217 45 -1183
rect 1613 -1217 1629 -1183
rect 29 -1233 1629 -1217
rect 1687 -1183 3287 -1145
rect 1687 -1217 1703 -1183
rect 3271 -1217 3287 -1183
rect 1687 -1233 3287 -1217
rect -3287 -1291 -1687 -1275
rect -3287 -1325 -3271 -1291
rect -1703 -1325 -1687 -1291
rect -3287 -1363 -1687 -1325
rect -1629 -1291 -29 -1275
rect -1629 -1325 -1613 -1291
rect -45 -1325 -29 -1291
rect -1629 -1363 -29 -1325
rect 29 -1291 1629 -1275
rect 29 -1325 45 -1291
rect 1613 -1325 1629 -1291
rect 29 -1363 1629 -1325
rect 1687 -1291 3287 -1275
rect 1687 -1325 1703 -1291
rect 3271 -1325 3287 -1291
rect 1687 -1363 3287 -1325
rect -3287 -1601 -1687 -1563
rect -3287 -1635 -3271 -1601
rect -1703 -1635 -1687 -1601
rect -3287 -1651 -1687 -1635
rect -1629 -1601 -29 -1563
rect -1629 -1635 -1613 -1601
rect -45 -1635 -29 -1601
rect -1629 -1651 -29 -1635
rect 29 -1601 1629 -1563
rect 29 -1635 45 -1601
rect 1613 -1635 1629 -1601
rect 29 -1651 1629 -1635
rect 1687 -1601 3287 -1563
rect 1687 -1635 1703 -1601
rect 3271 -1635 3287 -1601
rect 1687 -1651 3287 -1635
<< polycont >>
rect -3271 1601 -1703 1635
rect -1613 1601 -45 1635
rect 45 1601 1613 1635
rect 1703 1601 3271 1635
rect -3271 1291 -1703 1325
rect -1613 1291 -45 1325
rect 45 1291 1613 1325
rect 1703 1291 3271 1325
rect -3271 1183 -1703 1217
rect -1613 1183 -45 1217
rect 45 1183 1613 1217
rect 1703 1183 3271 1217
rect -3271 873 -1703 907
rect -1613 873 -45 907
rect 45 873 1613 907
rect 1703 873 3271 907
rect -3271 765 -1703 799
rect -1613 765 -45 799
rect 45 765 1613 799
rect 1703 765 3271 799
rect -3271 455 -1703 489
rect -1613 455 -45 489
rect 45 455 1613 489
rect 1703 455 3271 489
rect -3271 347 -1703 381
rect -1613 347 -45 381
rect 45 347 1613 381
rect 1703 347 3271 381
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect -3271 -381 -1703 -347
rect -1613 -381 -45 -347
rect 45 -381 1613 -347
rect 1703 -381 3271 -347
rect -3271 -489 -1703 -455
rect -1613 -489 -45 -455
rect 45 -489 1613 -455
rect 1703 -489 3271 -455
rect -3271 -799 -1703 -765
rect -1613 -799 -45 -765
rect 45 -799 1613 -765
rect 1703 -799 3271 -765
rect -3271 -907 -1703 -873
rect -1613 -907 -45 -873
rect 45 -907 1613 -873
rect 1703 -907 3271 -873
rect -3271 -1217 -1703 -1183
rect -1613 -1217 -45 -1183
rect 45 -1217 1613 -1183
rect 1703 -1217 3271 -1183
rect -3271 -1325 -1703 -1291
rect -1613 -1325 -45 -1291
rect 45 -1325 1613 -1291
rect 1703 -1325 3271 -1291
rect -3271 -1635 -1703 -1601
rect -1613 -1635 -45 -1601
rect 45 -1635 1613 -1601
rect 1703 -1635 3271 -1601
<< locali >>
rect -3447 1703 -3351 1737
rect 3351 1703 3447 1737
rect -3447 1641 -3413 1703
rect 3413 1641 3447 1703
rect -3287 1601 -3271 1635
rect -1703 1601 -1687 1635
rect -1629 1601 -1613 1635
rect -45 1601 -29 1635
rect 29 1601 45 1635
rect 1613 1601 1629 1635
rect 1687 1601 1703 1635
rect 3271 1601 3287 1635
rect -3333 1551 -3299 1567
rect -3333 1359 -3299 1375
rect -1675 1551 -1641 1567
rect -1675 1359 -1641 1375
rect -17 1551 17 1567
rect -17 1359 17 1375
rect 1641 1551 1675 1567
rect 1641 1359 1675 1375
rect 3299 1551 3333 1567
rect 3299 1359 3333 1375
rect -3287 1291 -3271 1325
rect -1703 1291 -1687 1325
rect -1629 1291 -1613 1325
rect -45 1291 -29 1325
rect 29 1291 45 1325
rect 1613 1291 1629 1325
rect 1687 1291 1703 1325
rect 3271 1291 3287 1325
rect -3287 1183 -3271 1217
rect -1703 1183 -1687 1217
rect -1629 1183 -1613 1217
rect -45 1183 -29 1217
rect 29 1183 45 1217
rect 1613 1183 1629 1217
rect 1687 1183 1703 1217
rect 3271 1183 3287 1217
rect -3333 1133 -3299 1149
rect -3333 941 -3299 957
rect -1675 1133 -1641 1149
rect -1675 941 -1641 957
rect -17 1133 17 1149
rect -17 941 17 957
rect 1641 1133 1675 1149
rect 1641 941 1675 957
rect 3299 1133 3333 1149
rect 3299 941 3333 957
rect -3287 873 -3271 907
rect -1703 873 -1687 907
rect -1629 873 -1613 907
rect -45 873 -29 907
rect 29 873 45 907
rect 1613 873 1629 907
rect 1687 873 1703 907
rect 3271 873 3287 907
rect -3287 765 -3271 799
rect -1703 765 -1687 799
rect -1629 765 -1613 799
rect -45 765 -29 799
rect 29 765 45 799
rect 1613 765 1629 799
rect 1687 765 1703 799
rect 3271 765 3287 799
rect -3333 715 -3299 731
rect -3333 523 -3299 539
rect -1675 715 -1641 731
rect -1675 523 -1641 539
rect -17 715 17 731
rect -17 523 17 539
rect 1641 715 1675 731
rect 1641 523 1675 539
rect 3299 715 3333 731
rect 3299 523 3333 539
rect -3287 455 -3271 489
rect -1703 455 -1687 489
rect -1629 455 -1613 489
rect -45 455 -29 489
rect 29 455 45 489
rect 1613 455 1629 489
rect 1687 455 1703 489
rect 3271 455 3287 489
rect -3287 347 -3271 381
rect -1703 347 -1687 381
rect -1629 347 -1613 381
rect -45 347 -29 381
rect 29 347 45 381
rect 1613 347 1629 381
rect 1687 347 1703 381
rect 3271 347 3287 381
rect -3333 297 -3299 313
rect -3333 105 -3299 121
rect -1675 297 -1641 313
rect -1675 105 -1641 121
rect -17 297 17 313
rect -17 105 17 121
rect 1641 297 1675 313
rect 1641 105 1675 121
rect 3299 297 3333 313
rect 3299 105 3333 121
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -1629 37 -1613 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1613 37 1629 71
rect 1687 37 1703 71
rect 3271 37 3287 71
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect -3333 -121 -3299 -105
rect -3333 -313 -3299 -297
rect -1675 -121 -1641 -105
rect -1675 -313 -1641 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 1641 -121 1675 -105
rect 1641 -313 1675 -297
rect 3299 -121 3333 -105
rect 3299 -313 3333 -297
rect -3287 -381 -3271 -347
rect -1703 -381 -1687 -347
rect -1629 -381 -1613 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 1613 -381 1629 -347
rect 1687 -381 1703 -347
rect 3271 -381 3287 -347
rect -3287 -489 -3271 -455
rect -1703 -489 -1687 -455
rect -1629 -489 -1613 -455
rect -45 -489 -29 -455
rect 29 -489 45 -455
rect 1613 -489 1629 -455
rect 1687 -489 1703 -455
rect 3271 -489 3287 -455
rect -3333 -539 -3299 -523
rect -3333 -731 -3299 -715
rect -1675 -539 -1641 -523
rect -1675 -731 -1641 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 1641 -539 1675 -523
rect 1641 -731 1675 -715
rect 3299 -539 3333 -523
rect 3299 -731 3333 -715
rect -3287 -799 -3271 -765
rect -1703 -799 -1687 -765
rect -1629 -799 -1613 -765
rect -45 -799 -29 -765
rect 29 -799 45 -765
rect 1613 -799 1629 -765
rect 1687 -799 1703 -765
rect 3271 -799 3287 -765
rect -3287 -907 -3271 -873
rect -1703 -907 -1687 -873
rect -1629 -907 -1613 -873
rect -45 -907 -29 -873
rect 29 -907 45 -873
rect 1613 -907 1629 -873
rect 1687 -907 1703 -873
rect 3271 -907 3287 -873
rect -3333 -957 -3299 -941
rect -3333 -1149 -3299 -1133
rect -1675 -957 -1641 -941
rect -1675 -1149 -1641 -1133
rect -17 -957 17 -941
rect -17 -1149 17 -1133
rect 1641 -957 1675 -941
rect 1641 -1149 1675 -1133
rect 3299 -957 3333 -941
rect 3299 -1149 3333 -1133
rect -3287 -1217 -3271 -1183
rect -1703 -1217 -1687 -1183
rect -1629 -1217 -1613 -1183
rect -45 -1217 -29 -1183
rect 29 -1217 45 -1183
rect 1613 -1217 1629 -1183
rect 1687 -1217 1703 -1183
rect 3271 -1217 3287 -1183
rect -3287 -1325 -3271 -1291
rect -1703 -1325 -1687 -1291
rect -1629 -1325 -1613 -1291
rect -45 -1325 -29 -1291
rect 29 -1325 45 -1291
rect 1613 -1325 1629 -1291
rect 1687 -1325 1703 -1291
rect 3271 -1325 3287 -1291
rect -3333 -1375 -3299 -1359
rect -3333 -1567 -3299 -1551
rect -1675 -1375 -1641 -1359
rect -1675 -1567 -1641 -1551
rect -17 -1375 17 -1359
rect -17 -1567 17 -1551
rect 1641 -1375 1675 -1359
rect 1641 -1567 1675 -1551
rect 3299 -1375 3333 -1359
rect 3299 -1567 3333 -1551
rect -3287 -1635 -3271 -1601
rect -1703 -1635 -1687 -1601
rect -1629 -1635 -1613 -1601
rect -45 -1635 -29 -1601
rect 29 -1635 45 -1601
rect 1613 -1635 1629 -1601
rect 1687 -1635 1703 -1601
rect 3271 -1635 3287 -1601
rect -3447 -1703 -3413 -1641
rect 3413 -1703 3447 -1641
rect -3447 -1737 -3351 -1703
rect 3351 -1737 3447 -1703
<< viali >>
rect -3271 1601 -1703 1635
rect -1613 1601 -45 1635
rect 45 1601 1613 1635
rect 1703 1601 3271 1635
rect -3333 1375 -3299 1551
rect -1675 1375 -1641 1551
rect -17 1375 17 1551
rect 1641 1375 1675 1551
rect 3299 1375 3333 1551
rect -3271 1291 -1703 1325
rect -1613 1291 -45 1325
rect 45 1291 1613 1325
rect 1703 1291 3271 1325
rect -3271 1183 -1703 1217
rect -1613 1183 -45 1217
rect 45 1183 1613 1217
rect 1703 1183 3271 1217
rect -3333 957 -3299 1133
rect -1675 957 -1641 1133
rect -17 957 17 1133
rect 1641 957 1675 1133
rect 3299 957 3333 1133
rect -3271 873 -1703 907
rect -1613 873 -45 907
rect 45 873 1613 907
rect 1703 873 3271 907
rect -3271 765 -1703 799
rect -1613 765 -45 799
rect 45 765 1613 799
rect 1703 765 3271 799
rect -3333 539 -3299 715
rect -1675 539 -1641 715
rect -17 539 17 715
rect 1641 539 1675 715
rect 3299 539 3333 715
rect -3271 455 -1703 489
rect -1613 455 -45 489
rect 45 455 1613 489
rect 1703 455 3271 489
rect -3271 347 -1703 381
rect -1613 347 -45 381
rect 45 347 1613 381
rect 1703 347 3271 381
rect -3333 121 -3299 297
rect -1675 121 -1641 297
rect -17 121 17 297
rect 1641 121 1675 297
rect 3299 121 3333 297
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect -3333 -297 -3299 -121
rect -1675 -297 -1641 -121
rect -17 -297 17 -121
rect 1641 -297 1675 -121
rect 3299 -297 3333 -121
rect -3271 -381 -1703 -347
rect -1613 -381 -45 -347
rect 45 -381 1613 -347
rect 1703 -381 3271 -347
rect -3271 -489 -1703 -455
rect -1613 -489 -45 -455
rect 45 -489 1613 -455
rect 1703 -489 3271 -455
rect -3333 -715 -3299 -539
rect -1675 -715 -1641 -539
rect -17 -715 17 -539
rect 1641 -715 1675 -539
rect 3299 -715 3333 -539
rect -3271 -799 -1703 -765
rect -1613 -799 -45 -765
rect 45 -799 1613 -765
rect 1703 -799 3271 -765
rect -3271 -907 -1703 -873
rect -1613 -907 -45 -873
rect 45 -907 1613 -873
rect 1703 -907 3271 -873
rect -3333 -1133 -3299 -957
rect -1675 -1133 -1641 -957
rect -17 -1133 17 -957
rect 1641 -1133 1675 -957
rect 3299 -1133 3333 -957
rect -3271 -1217 -1703 -1183
rect -1613 -1217 -45 -1183
rect 45 -1217 1613 -1183
rect 1703 -1217 3271 -1183
rect -3271 -1325 -1703 -1291
rect -1613 -1325 -45 -1291
rect 45 -1325 1613 -1291
rect 1703 -1325 3271 -1291
rect -3333 -1551 -3299 -1375
rect -1675 -1551 -1641 -1375
rect -17 -1551 17 -1375
rect 1641 -1551 1675 -1375
rect 3299 -1551 3333 -1375
rect -3271 -1635 -1703 -1601
rect -1613 -1635 -45 -1601
rect 45 -1635 1613 -1601
rect 1703 -1635 3271 -1601
<< metal1 >>
rect -3283 1635 -1691 1641
rect -3283 1601 -3271 1635
rect -1703 1601 -1691 1635
rect -3283 1595 -1691 1601
rect -1625 1635 -33 1641
rect -1625 1601 -1613 1635
rect -45 1601 -33 1635
rect -1625 1595 -33 1601
rect 33 1635 1625 1641
rect 33 1601 45 1635
rect 1613 1601 1625 1635
rect 33 1595 1625 1601
rect 1691 1635 3283 1641
rect 1691 1601 1703 1635
rect 3271 1601 3283 1635
rect 1691 1595 3283 1601
rect -3339 1551 -3293 1563
rect -3339 1375 -3333 1551
rect -3299 1375 -3293 1551
rect -3339 1363 -3293 1375
rect -1681 1551 -1635 1563
rect -1681 1375 -1675 1551
rect -1641 1375 -1635 1551
rect -1681 1363 -1635 1375
rect -23 1551 23 1563
rect -23 1375 -17 1551
rect 17 1375 23 1551
rect -23 1363 23 1375
rect 1635 1551 1681 1563
rect 1635 1375 1641 1551
rect 1675 1375 1681 1551
rect 1635 1363 1681 1375
rect 3293 1551 3339 1563
rect 3293 1375 3299 1551
rect 3333 1375 3339 1551
rect 3293 1363 3339 1375
rect -3283 1325 -1691 1331
rect -3283 1291 -3271 1325
rect -1703 1291 -1691 1325
rect -3283 1285 -1691 1291
rect -1625 1325 -33 1331
rect -1625 1291 -1613 1325
rect -45 1291 -33 1325
rect -1625 1285 -33 1291
rect 33 1325 1625 1331
rect 33 1291 45 1325
rect 1613 1291 1625 1325
rect 33 1285 1625 1291
rect 1691 1325 3283 1331
rect 1691 1291 1703 1325
rect 3271 1291 3283 1325
rect 1691 1285 3283 1291
rect -3283 1217 -1691 1223
rect -3283 1183 -3271 1217
rect -1703 1183 -1691 1217
rect -3283 1177 -1691 1183
rect -1625 1217 -33 1223
rect -1625 1183 -1613 1217
rect -45 1183 -33 1217
rect -1625 1177 -33 1183
rect 33 1217 1625 1223
rect 33 1183 45 1217
rect 1613 1183 1625 1217
rect 33 1177 1625 1183
rect 1691 1217 3283 1223
rect 1691 1183 1703 1217
rect 3271 1183 3283 1217
rect 1691 1177 3283 1183
rect -3339 1133 -3293 1145
rect -3339 957 -3333 1133
rect -3299 957 -3293 1133
rect -3339 945 -3293 957
rect -1681 1133 -1635 1145
rect -1681 957 -1675 1133
rect -1641 957 -1635 1133
rect -1681 945 -1635 957
rect -23 1133 23 1145
rect -23 957 -17 1133
rect 17 957 23 1133
rect -23 945 23 957
rect 1635 1133 1681 1145
rect 1635 957 1641 1133
rect 1675 957 1681 1133
rect 1635 945 1681 957
rect 3293 1133 3339 1145
rect 3293 957 3299 1133
rect 3333 957 3339 1133
rect 3293 945 3339 957
rect -3283 907 -1691 913
rect -3283 873 -3271 907
rect -1703 873 -1691 907
rect -3283 867 -1691 873
rect -1625 907 -33 913
rect -1625 873 -1613 907
rect -45 873 -33 907
rect -1625 867 -33 873
rect 33 907 1625 913
rect 33 873 45 907
rect 1613 873 1625 907
rect 33 867 1625 873
rect 1691 907 3283 913
rect 1691 873 1703 907
rect 3271 873 3283 907
rect 1691 867 3283 873
rect -3283 799 -1691 805
rect -3283 765 -3271 799
rect -1703 765 -1691 799
rect -3283 759 -1691 765
rect -1625 799 -33 805
rect -1625 765 -1613 799
rect -45 765 -33 799
rect -1625 759 -33 765
rect 33 799 1625 805
rect 33 765 45 799
rect 1613 765 1625 799
rect 33 759 1625 765
rect 1691 799 3283 805
rect 1691 765 1703 799
rect 3271 765 3283 799
rect 1691 759 3283 765
rect -3339 715 -3293 727
rect -3339 539 -3333 715
rect -3299 539 -3293 715
rect -3339 527 -3293 539
rect -1681 715 -1635 727
rect -1681 539 -1675 715
rect -1641 539 -1635 715
rect -1681 527 -1635 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 1635 715 1681 727
rect 1635 539 1641 715
rect 1675 539 1681 715
rect 1635 527 1681 539
rect 3293 715 3339 727
rect 3293 539 3299 715
rect 3333 539 3339 715
rect 3293 527 3339 539
rect -3283 489 -1691 495
rect -3283 455 -3271 489
rect -1703 455 -1691 489
rect -3283 449 -1691 455
rect -1625 489 -33 495
rect -1625 455 -1613 489
rect -45 455 -33 489
rect -1625 449 -33 455
rect 33 489 1625 495
rect 33 455 45 489
rect 1613 455 1625 489
rect 33 449 1625 455
rect 1691 489 3283 495
rect 1691 455 1703 489
rect 3271 455 3283 489
rect 1691 449 3283 455
rect -3283 381 -1691 387
rect -3283 347 -3271 381
rect -1703 347 -1691 381
rect -3283 341 -1691 347
rect -1625 381 -33 387
rect -1625 347 -1613 381
rect -45 347 -33 381
rect -1625 341 -33 347
rect 33 381 1625 387
rect 33 347 45 381
rect 1613 347 1625 381
rect 33 341 1625 347
rect 1691 381 3283 387
rect 1691 347 1703 381
rect 3271 347 3283 381
rect 1691 341 3283 347
rect -3339 297 -3293 309
rect -3339 121 -3333 297
rect -3299 121 -3293 297
rect -3339 109 -3293 121
rect -1681 297 -1635 309
rect -1681 121 -1675 297
rect -1641 121 -1635 297
rect -1681 109 -1635 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 1635 297 1681 309
rect 1635 121 1641 297
rect 1675 121 1681 297
rect 1635 109 1681 121
rect 3293 297 3339 309
rect 3293 121 3299 297
rect 3333 121 3339 297
rect 3293 109 3339 121
rect -3283 71 -1691 77
rect -3283 37 -3271 71
rect -1703 37 -1691 71
rect -3283 31 -1691 37
rect -1625 71 -33 77
rect -1625 37 -1613 71
rect -45 37 -33 71
rect -1625 31 -33 37
rect 33 71 1625 77
rect 33 37 45 71
rect 1613 37 1625 71
rect 33 31 1625 37
rect 1691 71 3283 77
rect 1691 37 1703 71
rect 3271 37 3283 71
rect 1691 31 3283 37
rect -3283 -37 -1691 -31
rect -3283 -71 -3271 -37
rect -1703 -71 -1691 -37
rect -3283 -77 -1691 -71
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect 1691 -37 3283 -31
rect 1691 -71 1703 -37
rect 3271 -71 3283 -37
rect 1691 -77 3283 -71
rect -3339 -121 -3293 -109
rect -3339 -297 -3333 -121
rect -3299 -297 -3293 -121
rect -3339 -309 -3293 -297
rect -1681 -121 -1635 -109
rect -1681 -297 -1675 -121
rect -1641 -297 -1635 -121
rect -1681 -309 -1635 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 1635 -121 1681 -109
rect 1635 -297 1641 -121
rect 1675 -297 1681 -121
rect 1635 -309 1681 -297
rect 3293 -121 3339 -109
rect 3293 -297 3299 -121
rect 3333 -297 3339 -121
rect 3293 -309 3339 -297
rect -3283 -347 -1691 -341
rect -3283 -381 -3271 -347
rect -1703 -381 -1691 -347
rect -3283 -387 -1691 -381
rect -1625 -347 -33 -341
rect -1625 -381 -1613 -347
rect -45 -381 -33 -347
rect -1625 -387 -33 -381
rect 33 -347 1625 -341
rect 33 -381 45 -347
rect 1613 -381 1625 -347
rect 33 -387 1625 -381
rect 1691 -347 3283 -341
rect 1691 -381 1703 -347
rect 3271 -381 3283 -347
rect 1691 -387 3283 -381
rect -3283 -455 -1691 -449
rect -3283 -489 -3271 -455
rect -1703 -489 -1691 -455
rect -3283 -495 -1691 -489
rect -1625 -455 -33 -449
rect -1625 -489 -1613 -455
rect -45 -489 -33 -455
rect -1625 -495 -33 -489
rect 33 -455 1625 -449
rect 33 -489 45 -455
rect 1613 -489 1625 -455
rect 33 -495 1625 -489
rect 1691 -455 3283 -449
rect 1691 -489 1703 -455
rect 3271 -489 3283 -455
rect 1691 -495 3283 -489
rect -3339 -539 -3293 -527
rect -3339 -715 -3333 -539
rect -3299 -715 -3293 -539
rect -3339 -727 -3293 -715
rect -1681 -539 -1635 -527
rect -1681 -715 -1675 -539
rect -1641 -715 -1635 -539
rect -1681 -727 -1635 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 1635 -539 1681 -527
rect 1635 -715 1641 -539
rect 1675 -715 1681 -539
rect 1635 -727 1681 -715
rect 3293 -539 3339 -527
rect 3293 -715 3299 -539
rect 3333 -715 3339 -539
rect 3293 -727 3339 -715
rect -3283 -765 -1691 -759
rect -3283 -799 -3271 -765
rect -1703 -799 -1691 -765
rect -3283 -805 -1691 -799
rect -1625 -765 -33 -759
rect -1625 -799 -1613 -765
rect -45 -799 -33 -765
rect -1625 -805 -33 -799
rect 33 -765 1625 -759
rect 33 -799 45 -765
rect 1613 -799 1625 -765
rect 33 -805 1625 -799
rect 1691 -765 3283 -759
rect 1691 -799 1703 -765
rect 3271 -799 3283 -765
rect 1691 -805 3283 -799
rect -3283 -873 -1691 -867
rect -3283 -907 -3271 -873
rect -1703 -907 -1691 -873
rect -3283 -913 -1691 -907
rect -1625 -873 -33 -867
rect -1625 -907 -1613 -873
rect -45 -907 -33 -873
rect -1625 -913 -33 -907
rect 33 -873 1625 -867
rect 33 -907 45 -873
rect 1613 -907 1625 -873
rect 33 -913 1625 -907
rect 1691 -873 3283 -867
rect 1691 -907 1703 -873
rect 3271 -907 3283 -873
rect 1691 -913 3283 -907
rect -3339 -957 -3293 -945
rect -3339 -1133 -3333 -957
rect -3299 -1133 -3293 -957
rect -3339 -1145 -3293 -1133
rect -1681 -957 -1635 -945
rect -1681 -1133 -1675 -957
rect -1641 -1133 -1635 -957
rect -1681 -1145 -1635 -1133
rect -23 -957 23 -945
rect -23 -1133 -17 -957
rect 17 -1133 23 -957
rect -23 -1145 23 -1133
rect 1635 -957 1681 -945
rect 1635 -1133 1641 -957
rect 1675 -1133 1681 -957
rect 1635 -1145 1681 -1133
rect 3293 -957 3339 -945
rect 3293 -1133 3299 -957
rect 3333 -1133 3339 -957
rect 3293 -1145 3339 -1133
rect -3283 -1183 -1691 -1177
rect -3283 -1217 -3271 -1183
rect -1703 -1217 -1691 -1183
rect -3283 -1223 -1691 -1217
rect -1625 -1183 -33 -1177
rect -1625 -1217 -1613 -1183
rect -45 -1217 -33 -1183
rect -1625 -1223 -33 -1217
rect 33 -1183 1625 -1177
rect 33 -1217 45 -1183
rect 1613 -1217 1625 -1183
rect 33 -1223 1625 -1217
rect 1691 -1183 3283 -1177
rect 1691 -1217 1703 -1183
rect 3271 -1217 3283 -1183
rect 1691 -1223 3283 -1217
rect -3283 -1291 -1691 -1285
rect -3283 -1325 -3271 -1291
rect -1703 -1325 -1691 -1291
rect -3283 -1331 -1691 -1325
rect -1625 -1291 -33 -1285
rect -1625 -1325 -1613 -1291
rect -45 -1325 -33 -1291
rect -1625 -1331 -33 -1325
rect 33 -1291 1625 -1285
rect 33 -1325 45 -1291
rect 1613 -1325 1625 -1291
rect 33 -1331 1625 -1325
rect 1691 -1291 3283 -1285
rect 1691 -1325 1703 -1291
rect 3271 -1325 3283 -1291
rect 1691 -1331 3283 -1325
rect -3339 -1375 -3293 -1363
rect -3339 -1551 -3333 -1375
rect -3299 -1551 -3293 -1375
rect -3339 -1563 -3293 -1551
rect -1681 -1375 -1635 -1363
rect -1681 -1551 -1675 -1375
rect -1641 -1551 -1635 -1375
rect -1681 -1563 -1635 -1551
rect -23 -1375 23 -1363
rect -23 -1551 -17 -1375
rect 17 -1551 23 -1375
rect -23 -1563 23 -1551
rect 1635 -1375 1681 -1363
rect 1635 -1551 1641 -1375
rect 1675 -1551 1681 -1375
rect 1635 -1563 1681 -1551
rect 3293 -1375 3339 -1363
rect 3293 -1551 3299 -1375
rect 3333 -1551 3339 -1375
rect 3293 -1563 3339 -1551
rect -3283 -1601 -1691 -1595
rect -3283 -1635 -3271 -1601
rect -1703 -1635 -1691 -1601
rect -3283 -1641 -1691 -1635
rect -1625 -1601 -33 -1595
rect -1625 -1635 -1613 -1601
rect -45 -1635 -33 -1601
rect -1625 -1641 -33 -1635
rect 33 -1601 1625 -1595
rect 33 -1635 45 -1601
rect 1613 -1635 1625 -1601
rect 33 -1641 1625 -1635
rect 1691 -1601 3283 -1595
rect 1691 -1635 1703 -1601
rect 3271 -1635 3283 -1601
rect 1691 -1641 3283 -1635
<< properties >>
string FIXED_BBOX -3430 -1720 3430 1720
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 8 m 8 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

../xspice/brownout_dig.out.spice